
module calc_DW_mult_tc_18 ( a, b, product, dw8_CLK );
  input [32:0] a;
  input [32:0] b;
  output [65:0] product;
  input dw8_CLK;
  wire   n6, n12, n15, n18, n21, n24, n27, n30, n33, n36, n39, n42, n44, n48,
         n50, n53, n55, n58, n61, n63, n66, n69, n71, n74, n77, n79, n82, n84,
         n86, n89, n91, n93, n95, n97, n99, n100, n102, n104, n105, n107, n109,
         n110, n112, n113, n114, n115, n116, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n149, n154, n155, n156, n157, n158, n160, n162, n163, n164,
         n165, n167, n169, n170, n172, n174, n175, n176, n177, n178, n179,
         n180, n182, n184, n185, n187, n189, n190, n191, n192, n197, n198,
         n199, n201, n205, n206, n207, n209, n211, n212, n214, n216, n218,
         n219, n220, n221, n222, n223, n224, n225, n227, n229, n230, n231,
         n232, n234, n237, n238, n239, n240, n242, n244, n245, n246, n247,
         n248, n249, n250, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n269, n271, n272,
         n274, n276, n277, n278, n280, n282, n283, n284, n285, n286, n288,
         n290, n291, n292, n293, n294, n296, n298, n299, n300, n301, n302,
         n304, n306, n308, n312, n319, n322, n324, n326, n327, n328, n329,
         n333, n335, n337, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1394, n1396, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1749, n1519, n1520, n1521, n1522,
         n1523, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748;
  assign n12 = a[3];
  assign n21 = a[5];
  assign n30 = a[7];
  assign n39 = a[9];
  assign n48 = a[11];
  assign n55 = a[13];
  assign n63 = a[15];
  assign n71 = a[17];
  assign n79 = a[19];
  assign n86 = a[21];
  assign n93 = a[23];
  assign n99 = a[25];
  assign n104 = a[27];
  assign n109 = a[29];
  assign n113 = a[32];
  assign n116 = b[0];
  assign n1358 = b[23];
  assign n1359 = b[22];
  assign n1360 = b[21];
  assign n1361 = b[20];
  assign n1362 = b[19];
  assign n1363 = b[18];
  assign n1364 = b[17];
  assign n1365 = b[16];
  assign n1366 = b[15];
  assign n1367 = b[14];
  assign n1368 = b[13];
  assign n1369 = b[12];
  assign n1370 = b[11];
  assign n1371 = b[10];
  assign n1372 = b[9];
  assign n1373 = b[8];
  assign n1374 = b[7];
  assign n1375 = b[6];
  assign n1376 = b[5];
  assign n1377 = b[4];
  assign n1378 = b[3];
  assign n1379 = b[2];
  assign n1380 = b[1];
  assign n1683 = dw8_CLK;

  CFA1X1 U97 ( .A(n383), .B(n1547), .CI(n356), .CO(n149), .S(product[30]) );
  CEO3X2 U346 ( .A(n359), .B(n341), .C(n357), .Z(n340) );
  CEO3X2 U347 ( .A(n361), .B(n1677), .C(n342), .Z(n341) );
  CEO3X2 U348 ( .A(n1676), .B(n363), .C(n344), .Z(n342) );
  CEO3X2 U349 ( .A(n347), .B(n346), .C(n365), .Z(n343) );
  CEO3X2 U350 ( .A(n1671), .B(n1675), .C(n1673), .Z(n344) );
  CEO3X2 U351 ( .A(n350), .B(n349), .C(n371), .Z(n345) );
  CEO3X2 U352 ( .A(n353), .B(n352), .C(n351), .Z(n346) );
  CEO3X2 U353 ( .A(n377), .B(n375), .C(n373), .Z(n347) );
  CEO3X2 U354 ( .A(n381), .B(n354), .C(n379), .Z(n348) );
  CEO3X2 U355 ( .A(n901), .B(n947), .C(n1031), .Z(n349) );
  CEO3X2 U356 ( .A(n863), .B(n923), .C(n1001), .Z(n350) );
  CEO3X2 U357 ( .A(n791), .B(n881), .C(n973), .Z(n351) );
  CEO3X2 U358 ( .A(n793), .B(n821), .C(n847), .Z(n352) );
  CEO3X2 U359 ( .A(n803), .B(n775), .C(n833), .Z(n353) );
  CFA1X1 U361 ( .A(n360), .B(n358), .CI(n385), .CO(n355), .S(n356) );
  CFA1X1 U362 ( .A(n364), .B(n387), .CI(n362), .CO(n357), .S(n358) );
  CFA1X1 U363 ( .A(n1674), .B(n389), .CI(n391), .CO(n359), .S(n360) );
  CFA1X1 U364 ( .A(n1668), .B(n1672), .CI(n1670), .CO(n361), .S(n362) );
  CFA1X1 U365 ( .A(n1664), .B(n1669), .CI(n1666), .CO(n363), .S(n364) );
  CFA1X1 U366 ( .A(n399), .B(n374), .CI(n376), .CO(n365), .S(n366) );
  CFA1X1 U367 ( .A(n382), .B(n378), .CI(n380), .CO(n367), .S(n368) );
  CFA1X1 U368 ( .A(n405), .B(n401), .CI(n403), .CO(n369), .S(n370) );
  CFA1X1 U369 ( .A(n948), .B(n407), .CI(n409), .CO(n371), .S(n372) );
  CFA1X1 U370 ( .A(n882), .B(n1002), .CI(n1032), .CO(n373), .S(n374) );
  CFA1X1 U371 ( .A(n864), .B(n974), .CI(n924), .CO(n375), .S(n376) );
  CFA1X1 U372 ( .A(n822), .B(n902), .CI(n848), .CO(n377), .S(n378) );
  CFA1X1 U373 ( .A(n794), .B(n834), .CI(n812), .CO(n379), .S(n380) );
  CFA1X1 U374 ( .A(n792), .B(n804), .CI(n798), .CO(n381), .S(n382) );
  CFA1X1 U375 ( .A(n388), .B(n386), .CI(n413), .CO(n383), .S(n384) );
  CFA1X1 U376 ( .A(n392), .B(n415), .CI(n390), .CO(n385), .S(n386) );
  CFA1X1 U377 ( .A(n1667), .B(n417), .CI(n1661), .CO(n387), .S(n388) );
  CFA1X1 U378 ( .A(n1663), .B(n1665), .CI(n1659), .CO(n389), .S(n390) );
  CFA1X1 U379 ( .A(n1662), .B(n1657), .CI(n1655), .CO(n391), .S(n392) );
  CFA1X1 U380 ( .A(n406), .B(n402), .CI(n404), .CO(n393), .S(n394) );
  CFA1X1 U381 ( .A(n427), .B(n408), .CI(n429), .CO(n395), .S(n396) );
  CFA1X1 U382 ( .A(n435), .B(n431), .CI(n433), .CO(n397), .S(n398) );
  CFA1X1 U383 ( .A(n949), .B(n410), .CI(n1033), .CO(n399), .S(n400) );
  CFA1X1 U384 ( .A(n865), .B(n975), .CI(n925), .CO(n401), .S(n402) );
  CFA1X1 U385 ( .A(n849), .B(n1003), .CI(n883), .CO(n403), .S(n404) );
  CFA1X1 U386 ( .A(n823), .B(n903), .CI(n795), .CO(n405), .S(n406) );
  CFA1X1 U387 ( .A(n805), .B(n835), .CI(n776), .CO(n407), .S(n408) );
  CHA1X1 U388 ( .A(n799), .B(n813), .CO(n409), .S(n410) );
  CFA1X1 U389 ( .A(n416), .B(n414), .CI(n439), .CO(n411), .S(n412) );
  CFA1X1 U390 ( .A(n1660), .B(n441), .CI(n418), .CO(n413), .S(n414) );
  CFA1X1 U391 ( .A(n1658), .B(n443), .CI(n445), .CO(n415), .S(n416) );
  CFA1X1 U392 ( .A(n1654), .B(n1656), .CI(n1653), .CO(n417), .S(n418) );
  CFA1X1 U393 ( .A(n428), .B(n449), .CI(n451), .CO(n419), .S(n420) );
  CFA1X1 U394 ( .A(n434), .B(n430), .CI(n432), .CO(n421), .S(n422) );
  CFA1X1 U395 ( .A(n455), .B(n436), .CI(n453), .CO(n423), .S(n424) );
  CFA1X1 U396 ( .A(n461), .B(n457), .CI(n459), .CO(n425), .S(n426) );
  CFA1X1 U397 ( .A(n904), .B(n1004), .CI(n926), .CO(n427), .S(n428) );
  CFA1X1 U398 ( .A(n884), .B(n976), .CI(n1034), .CO(n429), .S(n430) );
  CFA1X1 U399 ( .A(n836), .B(n950), .CI(n850), .CO(n431), .S(n432) );
  CFA1X1 U400 ( .A(n814), .B(n866), .CI(n824), .CO(n433), .S(n434) );
  CFA1X1 U401 ( .A(n796), .B(n806), .CI(n800), .CO(n435), .S(n436) );
  CFA1X1 U402 ( .A(n442), .B(n440), .CI(n465), .CO(n437), .S(n438) );
  CFA1X1 U403 ( .A(n446), .B(n467), .CI(n444), .CO(n439), .S(n440) );
  CFA1X1 U404 ( .A(n1647), .B(n469), .CI(n1652), .CO(n441), .S(n442) );
  CFA1X1 U405 ( .A(n1650), .B(n1651), .CI(n1645), .CO(n443), .S(n444) );
  CFA1X1 U406 ( .A(n1648), .B(n1643), .CI(n1649), .CO(n445), .S(n446) );
  CFA1X1 U407 ( .A(n460), .B(n456), .CI(n477), .CO(n447), .S(n448) );
  CFA1X1 U408 ( .A(n483), .B(n479), .CI(n481), .CO(n449), .S(n450) );
  CFA1X1 U409 ( .A(n927), .B(n485), .CI(n462), .CO(n451), .S(n452) );
  CFA1X1 U410 ( .A(n905), .B(n1005), .CI(n1035), .CO(n453), .S(n454) );
  CFA1X1 U411 ( .A(n851), .B(n977), .CI(n885), .CO(n455), .S(n456) );
  CFA1X1 U412 ( .A(n837), .B(n951), .CI(n801), .CO(n457), .S(n458) );
  CFA1X1 U413 ( .A(n815), .B(n867), .CI(n825), .CO(n459), .S(n460) );
  CHA1X1 U414 ( .A(n807), .B(n777), .CO(n461), .S(n462) );
  CFA1X1 U415 ( .A(n468), .B(n466), .CI(n489), .CO(n463), .S(n464) );
  CFA1X1 U416 ( .A(n493), .B(n491), .CI(n470), .CO(n465), .S(n466) );
  CFA1X1 U417 ( .A(n1641), .B(n1646), .CI(n1644), .CO(n467), .S(n468) );
  CFA1X1 U418 ( .A(n1637), .B(n1642), .CI(n1639), .CO(n469), .S(n470) );
  CFA1X1 U419 ( .A(n482), .B(n478), .CI(n480), .CO(n471), .S(n472) );
  CFA1X1 U420 ( .A(n503), .B(n484), .CI(n486), .CO(n473), .S(n474) );
  CFA1X1 U421 ( .A(n507), .B(n501), .CI(n505), .CO(n475), .S(n476) );
  CFA1X1 U422 ( .A(n928), .B(n509), .CI(n1006), .CO(n477), .S(n478) );
  CFA1X1 U423 ( .A(n886), .B(n978), .CI(n1036), .CO(n479), .S(n480) );
  CFA1X1 U424 ( .A(n838), .B(n952), .CI(n868), .CO(n481), .S(n482) );
  CFA1X1 U425 ( .A(n826), .B(n906), .CI(n852), .CO(n483), .S(n484) );
  CFA1X1 U426 ( .A(n802), .B(n816), .CI(n808), .CO(n485), .S(n486) );
  CFA1X1 U427 ( .A(n492), .B(n490), .CI(n513), .CO(n487), .S(n488) );
  CFA1X1 U428 ( .A(n517), .B(n515), .CI(n494), .CO(n489), .S(n490) );
  CFA1X1 U429 ( .A(n1635), .B(n1640), .CI(n1638), .CO(n491), .S(n492) );
  CFA1X1 U430 ( .A(n1631), .B(n1636), .CI(n1633), .CO(n493), .S(n494) );
  CFA1X1 U431 ( .A(n506), .B(n502), .CI(n504), .CO(n495), .S(n496) );
  CFA1X1 U432 ( .A(n527), .B(n508), .CI(n525), .CO(n497), .S(n498) );
  CFA1X1 U433 ( .A(n510), .B(n529), .CI(n531), .CO(n499), .S(n500) );
  CFA1X1 U434 ( .A(n929), .B(n1037), .CI(n953), .CO(n501), .S(n502) );
  CFA1X1 U435 ( .A(n809), .B(n979), .CI(n907), .CO(n503), .S(n504) );
  CFA1X1 U436 ( .A(n853), .B(n1007), .CI(n887), .CO(n505), .S(n506) );
  CFA1X1 U437 ( .A(n778), .B(n869), .CI(n839), .CO(n507), .S(n508) );
  CHA1X1 U438 ( .A(n817), .B(n827), .CO(n509), .S(n510) );
  CFA1X1 U439 ( .A(n516), .B(n514), .CI(n535), .CO(n511), .S(n512) );
  CFA1X1 U441 ( .A(n1626), .B(n1634), .CI(n1632), .CO(n515), .S(n516) );
  CFA1X1 U443 ( .A(n530), .B(n545), .CI(n528), .CO(n519), .S(n520) );
  CFA1X1 U444 ( .A(n549), .B(n532), .CI(n547), .CO(n521), .S(n522) );
  CFA1X1 U445 ( .A(n930), .B(n551), .CI(n553), .CO(n523), .S(n524) );
  CFA1X1 U446 ( .A(n908), .B(n980), .CI(n1038), .CO(n525), .S(n526) );
  CFA1X1 U447 ( .A(n854), .B(n1008), .CI(n888), .CO(n527), .S(n528) );
  CFA1X1 U448 ( .A(n840), .B(n954), .CI(n870), .CO(n529), .S(n530) );
  CFA1X1 U449 ( .A(n810), .B(n828), .CI(n818), .CO(n531), .S(n532) );
  CFA1X1 U450 ( .A(n538), .B(n536), .CI(n557), .CO(n533), .S(n534) );
  CFA1X1 U451 ( .A(n1625), .B(n559), .CI(n1627), .CO(n535), .S(n536) );
  CFA1X1 U452 ( .A(n1620), .B(n1622), .CI(n1623), .CO(n537), .S(n538) );
  CFA1X1 U453 ( .A(n548), .B(n565), .CI(n546), .CO(n539), .S(n540) );
  CFA1X1 U454 ( .A(n567), .B(n550), .CI(n552), .CO(n541), .S(n542) );
  CFA1X1 U455 ( .A(n573), .B(n569), .CI(n571), .CO(n543), .S(n544) );
  CFA1X1 U456 ( .A(n931), .B(n554), .CI(n1039), .CO(n545), .S(n546) );
  CFA1X1 U457 ( .A(n819), .B(n981), .CI(n909), .CO(n547), .S(n548) );
  CFA1X1 U458 ( .A(n855), .B(n1009), .CI(n889), .CO(n549), .S(n550) );
  CFA1X1 U459 ( .A(n841), .B(n955), .CI(n871), .CO(n551), .S(n552) );
  CHA1X1 U460 ( .A(n779), .B(n829), .CO(n553), .S(n554) );
  CFA1X1 U461 ( .A(n560), .B(n558), .CI(n577), .CO(n555), .S(n556) );
  CFA1X1 U462 ( .A(n1619), .B(n579), .CI(n1621), .CO(n557), .S(n558) );
  CFA1X1 U463 ( .A(n1615), .B(n1617), .CI(n1618), .CO(n559), .S(n560) );
  CFA1X1 U464 ( .A(n570), .B(n585), .CI(n568), .CO(n561), .S(n562) );
  CFA1X1 U465 ( .A(n587), .B(n572), .CI(n574), .CO(n563), .S(n564) );
  CFA1X1 U466 ( .A(n593), .B(n589), .CI(n591), .CO(n565), .S(n566) );
  CFA1X1 U467 ( .A(n910), .B(n1040), .CI(n956), .CO(n567), .S(n568) );
  CFA1X1 U468 ( .A(n872), .B(n1010), .CI(n932), .CO(n569), .S(n570) );
  CFA1X1 U469 ( .A(n856), .B(n982), .CI(n890), .CO(n571), .S(n572) );
  CFA1X1 U470 ( .A(n820), .B(n842), .CI(n830), .CO(n573), .S(n574) );
  CFA1X1 U471 ( .A(n580), .B(n578), .CI(n597), .CO(n575), .S(n576) );
  CFA1X1 U472 ( .A(n1614), .B(n599), .CI(n1616), .CO(n577), .S(n578) );
  CFA1X1 U473 ( .A(n1610), .B(n1612), .CI(n1613), .CO(n579), .S(n580) );
  CFA1X1 U474 ( .A(n605), .B(n588), .CI(n590), .CO(n581), .S(n582) );
  CFA1X1 U475 ( .A(n609), .B(n592), .CI(n607), .CO(n583), .S(n584) );
  CFA1X1 U476 ( .A(n933), .B(n611), .CI(n594), .CO(n585), .S(n586) );
  CFA1X1 U477 ( .A(n911), .B(n1011), .CI(n1041), .CO(n587), .S(n588) );
  CFA1X1 U478 ( .A(n857), .B(n983), .CI(n891), .CO(n589), .S(n590) );
  CFA1X1 U479 ( .A(n843), .B(n957), .CI(n873), .CO(n591), .S(n592) );
  CHA1X1 U480 ( .A(n780), .B(n831), .CO(n593), .S(n594) );
  CFA1X1 U481 ( .A(n600), .B(n598), .CI(n615), .CO(n595), .S(n596) );
  CFA1X1 U482 ( .A(n1609), .B(n617), .CI(n1611), .CO(n597), .S(n598) );
  CFA1X1 U483 ( .A(n1608), .B(n1607), .CI(n1605), .CO(n599), .S(n600) );
  CFA1X1 U484 ( .A(n612), .B(n608), .CI(n610), .CO(n601), .S(n602) );
  CFA1X1 U485 ( .A(n627), .B(n623), .CI(n625), .CO(n603), .S(n604) );
  CFA1X1 U486 ( .A(n912), .B(n629), .CI(n958), .CO(n605), .S(n606) );
  CFA1X1 U487 ( .A(n892), .B(n1012), .CI(n1042), .CO(n607), .S(n608) );
  CFA1X1 U488 ( .A(n874), .B(n984), .CI(n934), .CO(n609), .S(n610) );
  CFA1X1 U489 ( .A(n832), .B(n858), .CI(n844), .CO(n611), .S(n612) );
  CFA1X1 U490 ( .A(n618), .B(n616), .CI(n633), .CO(n613), .S(n614) );
  CFA1X1 U491 ( .A(n1604), .B(n1602), .CI(n1606), .CO(n615), .S(n616) );
  CFA1X1 U492 ( .A(n1603), .B(n1600), .CI(n1598), .CO(n617), .S(n618) );
  CFA1X1 U493 ( .A(n643), .B(n626), .CI(n628), .CO(n619), .S(n620) );
  CFA1X1 U494 ( .A(n630), .B(n641), .CI(n645), .CO(n621), .S(n622) );
  CFA1X1 U495 ( .A(n935), .B(n1043), .CI(n959), .CO(n623), .S(n624) );
  CFA1X1 U496 ( .A(n845), .B(n1013), .CI(n913), .CO(n625), .S(n626) );
  CFA1X1 U497 ( .A(n859), .B(n985), .CI(n893), .CO(n627), .S(n628) );
  CHA1X1 U498 ( .A(n781), .B(n875), .CO(n629), .S(n630) );
  CFA1X1 U499 ( .A(n1601), .B(n634), .CI(n649), .CO(n631), .S(n632) );
  CFA1X1 U500 ( .A(n1597), .B(n1596), .CI(n1599), .CO(n633), .S(n634) );
  CFA1X1 U501 ( .A(n642), .B(n653), .CI(n655), .CO(n635), .S(n636) );
  CFA1X1 U502 ( .A(n657), .B(n644), .CI(n646), .CO(n637), .S(n638) );
  CFA1X1 U503 ( .A(n936), .B(n659), .CI(n661), .CO(n639), .S(n640) );
  CFA1X1 U504 ( .A(n914), .B(n1014), .CI(n960), .CO(n641), .S(n642) );
  CFA1X1 U505 ( .A(n894), .B(n986), .CI(n1044), .CO(n643), .S(n644) );
  CFA1X1 U506 ( .A(n846), .B(n876), .CI(n860), .CO(n645), .S(n646) );
  CFA1X1 U507 ( .A(n1595), .B(n650), .CI(n1593), .CO(n647), .S(n648) );
  CFA1X1 U508 ( .A(n1589), .B(n1591), .CI(n1594), .CO(n649), .S(n650) );
  CFA1X1 U509 ( .A(n660), .B(n656), .CI(n658), .CO(n651), .S(n652) );
  CFA1X1 U510 ( .A(n675), .B(n673), .CI(n671), .CO(n653), .S(n654) );
  CFA1X1 U511 ( .A(n895), .B(n662), .CI(n1045), .CO(n655), .S(n656) );
  CFA1X1 U512 ( .A(n861), .B(n1015), .CI(n961), .CO(n657), .S(n658) );
  CFA1X1 U513 ( .A(n877), .B(n987), .CI(n937), .CO(n659), .S(n660) );
  CHA1X1 U514 ( .A(n782), .B(n915), .CO(n661), .S(n662) );
  CFA1X1 U515 ( .A(n1590), .B(n1592), .CI(n1588), .CO(n663), .S(n664) );
  CFA1X1 U516 ( .A(n683), .B(n681), .CI(n670), .CO(n665), .S(n666) );
  CFA1X1 U517 ( .A(n676), .B(n672), .CI(n674), .CO(n667), .S(n668) );
  CFA1X1 U518 ( .A(n689), .B(n685), .CI(n687), .CO(n669), .S(n670) );
  CFA1X1 U519 ( .A(n938), .B(n1046), .CI(n962), .CO(n671), .S(n672) );
  CFA1X1 U520 ( .A(n916), .B(n1016), .CI(n988), .CO(n673), .S(n674) );
  CFA1X1 U521 ( .A(n862), .B(n896), .CI(n878), .CO(n675), .S(n676) );
  CFA1X1 U522 ( .A(n1586), .B(n1587), .CI(n1585), .CO(n677), .S(n678) );
  CFA1X1 U523 ( .A(n697), .B(n684), .CI(n695), .CO(n679), .S(n680) );
  CFA1X1 U524 ( .A(n699), .B(n686), .CI(n688), .CO(n681), .S(n682) );
  CFA1X1 U525 ( .A(n917), .B(n701), .CI(n690), .CO(n683), .S(n684) );
  CFA1X1 U526 ( .A(n897), .B(n989), .CI(n1047), .CO(n685), .S(n686) );
  CFA1X1 U527 ( .A(n879), .B(n1017), .CI(n963), .CO(n687), .S(n688) );
  CHA1X1 U528 ( .A(n783), .B(n939), .CO(n689), .S(n690) );
  CFA1X1 U529 ( .A(n1583), .B(n1584), .CI(n1582), .CO(n691), .S(n692) );
  CFA1X1 U530 ( .A(n700), .B(n707), .CI(n698), .CO(n693), .S(n694) );
  CFA1X1 U531 ( .A(n709), .B(n702), .CI(n711), .CO(n695), .S(n696) );
  CFA1X1 U532 ( .A(n964), .B(n713), .CI(n1048), .CO(n697), .S(n698) );
  CFA1X1 U533 ( .A(n940), .B(n990), .CI(n1018), .CO(n699), .S(n700) );
  CFA1X1 U534 ( .A(n880), .B(n918), .CI(n898), .CO(n701), .S(n702) );
  CFA1X1 U535 ( .A(n1580), .B(n1581), .CI(n1579), .CO(n703), .S(n704) );
  CFA1X1 U536 ( .A(n712), .B(n719), .CI(n710), .CO(n705), .S(n706) );
  CFA1X1 U537 ( .A(n714), .B(n721), .CI(n723), .CO(n707), .S(n708) );
  CFA1X1 U538 ( .A(n919), .B(n965), .CI(n941), .CO(n709), .S(n710) );
  CFA1X1 U539 ( .A(n899), .B(n991), .CI(n1049), .CO(n711), .S(n712) );
  CHA1X1 U540 ( .A(n784), .B(n1019), .CO(n713), .S(n714) );
  CFA1X1 U541 ( .A(n1576), .B(n1578), .CI(n1577), .CO(n715), .S(n716) );
  CFA1X1 U542 ( .A(n724), .B(n729), .CI(n722), .CO(n717), .S(n718) );
  CFA1X1 U543 ( .A(n1050), .B(n731), .CI(n733), .CO(n719), .S(n720) );
  CFA1X1 U544 ( .A(n966), .B(n1020), .CI(n992), .CO(n721), .S(n722) );
  CFA1X1 U545 ( .A(n900), .B(n942), .CI(n920), .CO(n723), .S(n724) );
  CFA1X1 U546 ( .A(n1574), .B(n1575), .CI(n1573), .CO(n725), .S(n726) );
  CFA1X1 U547 ( .A(n741), .B(n732), .CI(n739), .CO(n727), .S(n728) );
  CFA1X1 U548 ( .A(n943), .B(n734), .CI(n967), .CO(n729), .S(n730) );
  CFA1X1 U549 ( .A(n921), .B(n993), .CI(n1051), .CO(n731), .S(n732) );
  CHA1X1 U550 ( .A(n785), .B(n1021), .CO(n733), .S(n734) );
  CFA1X1 U551 ( .A(n1571), .B(n1572), .CI(n1568), .CO(n735), .S(n736) );
  CFA1X1 U552 ( .A(n749), .B(n742), .CI(n747), .CO(n737), .S(n738) );
  CFA1X1 U553 ( .A(n1052), .B(n1022), .CI(n994), .CO(n739), .S(n740) );
  CFA1X1 U554 ( .A(n922), .B(n968), .CI(n944), .CO(n741), .S(n742) );
  CFA1X1 U555 ( .A(n753), .B(n746), .CI(n748), .CO(n743), .S(n744) );
  CFA1X1 U556 ( .A(n969), .B(n755), .CI(n750), .CO(n745), .S(n746) );
  CFA1X1 U557 ( .A(n945), .B(n995), .CI(n1053), .CO(n747), .S(n748) );
  CHA1X1 U558 ( .A(n786), .B(n1023), .CO(n749), .S(n750) );
  CFA1X1 U559 ( .A(n759), .B(n754), .CI(n756), .CO(n751), .S(n752) );
  CFA1X1 U560 ( .A(n1024), .B(n761), .CI(n996), .CO(n753), .S(n754) );
  CFA1X1 U561 ( .A(n946), .B(n1054), .CI(n970), .CO(n755), .S(n756) );
  CFA1X1 U562 ( .A(n762), .B(n760), .CI(n765), .CO(n757), .S(n758) );
  CFA1X1 U563 ( .A(n971), .B(n997), .CI(n1055), .CO(n759), .S(n760) );
  CHA1X1 U564 ( .A(n787), .B(n1025), .CO(n761), .S(n762) );
  CFA1X1 U565 ( .A(n998), .B(n766), .CI(n769), .CO(n763), .S(n764) );
  CFA1X1 U566 ( .A(n972), .B(n1026), .CI(n1056), .CO(n765), .S(n766) );
  CFA1X1 U567 ( .A(n1027), .B(n770), .CI(n999), .CO(n767), .S(n768) );
  CHA1X1 U568 ( .A(n1057), .B(n788), .CO(n769), .S(n770) );
  CFA1X1 U569 ( .A(n1000), .B(n1028), .CI(n1058), .CO(n771), .S(n772) );
  CHA1X1 U570 ( .A(n1059), .B(n1029), .CO(n773), .S(n774) );
  COND2X1 U571 ( .A(n115), .B(n1407), .C(n114), .D(n1064), .Z(n775) );
  COND2X1 U572 ( .A(n1063), .B(n115), .C(n114), .D(n1062), .Z(n791) );
  COND2X1 U578 ( .A(n112), .B(n1066), .C(n110), .D(n1065), .Z(n793) );
  COND2X1 U580 ( .A(n1068), .B(n112), .C(n110), .D(n1067), .Z(n795) );
  COND2X1 U589 ( .A(n107), .B(n1072), .C(n105), .D(n1071), .Z(n798) );
  COND2X1 U592 ( .A(n1075), .B(n107), .C(n105), .D(n1074), .Z(n801) );
  COND2X1 U601 ( .A(n102), .B(n1410), .C(n100), .D(n1085), .Z(n778) );
  COND2X1 U602 ( .A(n102), .B(n1078), .C(n100), .D(n1077), .Z(n803) );
  COND2X1 U603 ( .A(n102), .B(n1079), .C(n100), .D(n1078), .Z(n804) );
  COND2X1 U605 ( .A(n102), .B(n1081), .C(n100), .D(n1080), .Z(n806) );
  COND2X1 U608 ( .A(n1084), .B(n102), .C(n100), .D(n1083), .Z(n809) );
  COND2X1 U619 ( .A(n97), .B(n1411), .C(n95), .D(n1096), .Z(n779) );
  COND2X1 U620 ( .A(n97), .B(n1087), .C(n1086), .D(n95), .Z(n811) );
  COND2X1 U623 ( .A(n97), .B(n1090), .C(n1089), .D(n95), .Z(n814) );
  COND2X1 U624 ( .A(n97), .B(n1091), .C(n1090), .D(n95), .Z(n815) );
  COND2X1 U625 ( .A(n97), .B(n1092), .C(n1091), .D(n95), .Z(n816) );
  COND2X1 U626 ( .A(n97), .B(n1093), .C(n1092), .D(n95), .Z(n817) );
  COND2X1 U628 ( .A(n1095), .B(n97), .C(n95), .D(n1094), .Z(n819) );
  COND2X1 U641 ( .A(n91), .B(n1412), .C(n89), .D(n1109), .Z(n780) );
  COND2X1 U642 ( .A(n91), .B(n1098), .C(n1097), .D(n89), .Z(n821) );
  COND2X1 U643 ( .A(n91), .B(n1099), .C(n1098), .D(n89), .Z(n822) );
  COND2X1 U644 ( .A(n91), .B(n1100), .C(n1099), .D(n89), .Z(n823) );
  COND2X1 U645 ( .A(n91), .B(n1101), .C(n1100), .D(n89), .Z(n824) );
  COND2X1 U646 ( .A(n91), .B(n1102), .C(n1101), .D(n89), .Z(n825) );
  COND2X1 U647 ( .A(n91), .B(n1103), .C(n1102), .D(n89), .Z(n826) );
  COND2X1 U648 ( .A(n91), .B(n1104), .C(n1103), .D(n89), .Z(n827) );
  COND2X1 U649 ( .A(n91), .B(n1105), .C(n1104), .D(n89), .Z(n828) );
  COND2X1 U650 ( .A(n91), .B(n1106), .C(n1105), .D(n89), .Z(n829) );
  COND2X1 U652 ( .A(n1108), .B(n91), .C(n1107), .D(n89), .Z(n831) );
  COND2X1 U667 ( .A(n84), .B(n1413), .C(n82), .D(n1124), .Z(n781) );
  COND2X1 U668 ( .A(n84), .B(n1111), .C(n1110), .D(n82), .Z(n833) );
  COND2X1 U671 ( .A(n84), .B(n1114), .C(n1113), .D(n82), .Z(n836) );
  COND2X1 U672 ( .A(n84), .B(n1115), .C(n1114), .D(n82), .Z(n837) );
  COND2X1 U673 ( .A(n84), .B(n1116), .C(n1115), .D(n82), .Z(n838) );
  COND2X1 U674 ( .A(n84), .B(n1117), .C(n1116), .D(n82), .Z(n839) );
  COND2X1 U675 ( .A(n84), .B(n1118), .C(n1117), .D(n82), .Z(n840) );
  COND2X1 U676 ( .A(n84), .B(n1119), .C(n1118), .D(n82), .Z(n841) );
  COND2X1 U677 ( .A(n84), .B(n1120), .C(n1119), .D(n82), .Z(n842) );
  COND2X1 U678 ( .A(n84), .B(n1121), .C(n1120), .D(n82), .Z(n843) );
  COND2X1 U680 ( .A(n1123), .B(n84), .C(n1122), .D(n82), .Z(n845) );
  CND2IX1 U696 ( .B(n1748), .A(n1701), .Z(n1124) );
  COND2X1 U697 ( .A(n77), .B(n1414), .C(n74), .D(n1141), .Z(n782) );
  COND2X1 U698 ( .A(n77), .B(n1126), .C(n1125), .D(n74), .Z(n847) );
  COND2X1 U699 ( .A(n77), .B(n1127), .C(n1126), .D(n74), .Z(n848) );
  COND2X1 U700 ( .A(n77), .B(n1128), .C(n1127), .D(n74), .Z(n849) );
  COND2X1 U701 ( .A(n77), .B(n1129), .C(n1128), .D(n74), .Z(n850) );
  COND2X1 U702 ( .A(n77), .B(n1130), .C(n1129), .D(n74), .Z(n851) );
  COND2X1 U703 ( .A(n77), .B(n1131), .C(n1130), .D(n74), .Z(n852) );
  COND2X1 U704 ( .A(n77), .B(n1132), .C(n1131), .D(n74), .Z(n853) );
  COND2X1 U705 ( .A(n77), .B(n1133), .C(n1132), .D(n74), .Z(n854) );
  COND2X1 U706 ( .A(n77), .B(n1134), .C(n1133), .D(n74), .Z(n855) );
  COND2X1 U707 ( .A(n77), .B(n1135), .C(n1134), .D(n74), .Z(n856) );
  COND2X1 U708 ( .A(n77), .B(n1136), .C(n1135), .D(n74), .Z(n857) );
  COND2X1 U709 ( .A(n77), .B(n1137), .C(n1136), .D(n74), .Z(n858) );
  COND2X1 U710 ( .A(n77), .B(n1138), .C(n1137), .D(n74), .Z(n859) );
  COND2X1 U711 ( .A(n77), .B(n1139), .C(n1138), .D(n74), .Z(n860) );
  COND2X1 U712 ( .A(n1140), .B(n77), .C(n1139), .D(n74), .Z(n861) );
  COND2X1 U731 ( .A(n69), .B(n1415), .C(n1160), .D(n66), .Z(n783) );
  COND2X1 U732 ( .A(n69), .B(n1143), .C(n1142), .D(n66), .Z(n863) );
  COND2X1 U733 ( .A(n69), .B(n1144), .C(n1143), .D(n66), .Z(n864) );
  COND2X1 U734 ( .A(n69), .B(n1145), .C(n1144), .D(n66), .Z(n865) );
  COND2X1 U735 ( .A(n69), .B(n1146), .C(n1145), .D(n66), .Z(n866) );
  COND2X1 U736 ( .A(n69), .B(n1147), .C(n1146), .D(n66), .Z(n867) );
  COND2X1 U737 ( .A(n69), .B(n1148), .C(n1147), .D(n66), .Z(n868) );
  COND2X1 U738 ( .A(n69), .B(n1149), .C(n1148), .D(n66), .Z(n869) );
  COND2X1 U739 ( .A(n69), .B(n1150), .C(n1149), .D(n66), .Z(n870) );
  COND2X1 U740 ( .A(n69), .B(n1151), .C(n1150), .D(n66), .Z(n871) );
  COND2X1 U741 ( .A(n69), .B(n1152), .C(n1151), .D(n66), .Z(n872) );
  COND2X1 U742 ( .A(n69), .B(n1153), .C(n1152), .D(n66), .Z(n873) );
  COND2X1 U743 ( .A(n69), .B(n1154), .C(n1153), .D(n66), .Z(n874) );
  COND2X1 U744 ( .A(n69), .B(n1155), .C(n1154), .D(n66), .Z(n875) );
  COND2X1 U746 ( .A(n69), .B(n1157), .C(n1156), .D(n66), .Z(n877) );
  COND2X1 U748 ( .A(n69), .B(n1159), .C(n1158), .D(n66), .Z(n879) );
  CND2IX1 U768 ( .B(n1748), .A(n1699), .Z(n1160) );
  COND2X1 U769 ( .A(n61), .B(n1746), .C(n1181), .D(n58), .Z(n784) );
  COND2X1 U770 ( .A(n61), .B(n1162), .C(n1161), .D(n58), .Z(n881) );
  COND2X1 U771 ( .A(n61), .B(n1163), .C(n1162), .D(n58), .Z(n882) );
  COND2X1 U772 ( .A(n61), .B(n1164), .C(n1163), .D(n58), .Z(n883) );
  COND2X1 U773 ( .A(n61), .B(n1165), .C(n1164), .D(n58), .Z(n884) );
  COND2X1 U774 ( .A(n61), .B(n1166), .C(n1165), .D(n58), .Z(n885) );
  COND2X1 U775 ( .A(n61), .B(n1167), .C(n1166), .D(n58), .Z(n886) );
  COND2X1 U776 ( .A(n61), .B(n1168), .C(n1167), .D(n58), .Z(n887) );
  COND2X1 U777 ( .A(n61), .B(n1169), .C(n1168), .D(n58), .Z(n888) );
  COND2X1 U778 ( .A(n61), .B(n1170), .C(n1169), .D(n58), .Z(n889) );
  COND2X1 U779 ( .A(n61), .B(n1171), .C(n1170), .D(n58), .Z(n890) );
  COND2X1 U780 ( .A(n61), .B(n1172), .C(n1171), .D(n58), .Z(n891) );
  COND2X1 U781 ( .A(n61), .B(n1173), .C(n1172), .D(n58), .Z(n892) );
  COND2X1 U782 ( .A(n61), .B(n1174), .C(n1173), .D(n58), .Z(n893) );
  COND2X1 U783 ( .A(n61), .B(n1175), .C(n1174), .D(n58), .Z(n894) );
  COND2X1 U784 ( .A(n61), .B(n1176), .C(n1175), .D(n58), .Z(n895) );
  COND2X1 U785 ( .A(n61), .B(n1177), .C(n1176), .D(n58), .Z(n896) );
  COND2X1 U786 ( .A(n61), .B(n1178), .C(n1177), .D(n58), .Z(n897) );
  COND2X1 U787 ( .A(n61), .B(n1179), .C(n1178), .D(n58), .Z(n898) );
  COND2X1 U788 ( .A(n61), .B(n1180), .C(n1179), .D(n58), .Z(n899) );
  CND2IX1 U810 ( .B(n1748), .A(n1745), .Z(n1181) );
  COND2X1 U811 ( .A(n53), .B(n1743), .C(n1204), .D(n50), .Z(n785) );
  COND2X1 U812 ( .A(n53), .B(n1183), .C(n1182), .D(n50), .Z(n901) );
  COND2X1 U813 ( .A(n53), .B(n1184), .C(n1183), .D(n50), .Z(n902) );
  COND2X1 U814 ( .A(n53), .B(n1185), .C(n1184), .D(n50), .Z(n903) );
  COND2X1 U815 ( .A(n53), .B(n1186), .C(n1185), .D(n50), .Z(n904) );
  COND2X1 U816 ( .A(n53), .B(n1187), .C(n1186), .D(n50), .Z(n905) );
  COND2X1 U817 ( .A(n53), .B(n1188), .C(n1187), .D(n50), .Z(n906) );
  COND2X1 U818 ( .A(n53), .B(n1189), .C(n1188), .D(n50), .Z(n907) );
  COND2X1 U819 ( .A(n53), .B(n1190), .C(n1189), .D(n50), .Z(n908) );
  COND2X1 U820 ( .A(n53), .B(n1191), .C(n1190), .D(n50), .Z(n909) );
  COND2X1 U821 ( .A(n53), .B(n1192), .C(n1191), .D(n50), .Z(n910) );
  COND2X1 U822 ( .A(n53), .B(n1193), .C(n1192), .D(n50), .Z(n911) );
  COND2X1 U823 ( .A(n53), .B(n1194), .C(n1193), .D(n50), .Z(n912) );
  COND2X1 U824 ( .A(n53), .B(n1195), .C(n1194), .D(n50), .Z(n913) );
  COND2X1 U825 ( .A(n53), .B(n1196), .C(n1195), .D(n50), .Z(n914) );
  COND2X1 U826 ( .A(n53), .B(n1197), .C(n1196), .D(n50), .Z(n915) );
  COND2X1 U827 ( .A(n53), .B(n1198), .C(n1197), .D(n50), .Z(n916) );
  COND2X1 U828 ( .A(n53), .B(n1199), .C(n1198), .D(n50), .Z(n917) );
  COND2X1 U829 ( .A(n53), .B(n1200), .C(n1199), .D(n50), .Z(n918) );
  COND2X1 U830 ( .A(n53), .B(n1201), .C(n1200), .D(n50), .Z(n919) );
  COND2X1 U831 ( .A(n53), .B(n1202), .C(n1201), .D(n50), .Z(n920) );
  COND2X1 U832 ( .A(n53), .B(n1203), .C(n1202), .D(n50), .Z(n921) );
  CND2IX1 U856 ( .B(n1748), .A(n1742), .Z(n1204) );
  COND2X1 U857 ( .A(n44), .B(n1738), .C(n1229), .D(n42), .Z(n786) );
  COND2X1 U858 ( .A(n44), .B(n1206), .C(n1205), .D(n42), .Z(n923) );
  COND2X1 U859 ( .A(n44), .B(n1207), .C(n1206), .D(n42), .Z(n924) );
  COND2X1 U860 ( .A(n44), .B(n1208), .C(n1207), .D(n42), .Z(n925) );
  COND2X1 U861 ( .A(n44), .B(n1209), .C(n1208), .D(n42), .Z(n926) );
  COND2X1 U862 ( .A(n44), .B(n1210), .C(n1209), .D(n42), .Z(n927) );
  COND2X1 U863 ( .A(n44), .B(n1211), .C(n1210), .D(n42), .Z(n928) );
  COND2X1 U864 ( .A(n44), .B(n1212), .C(n1211), .D(n42), .Z(n929) );
  COND2X1 U865 ( .A(n44), .B(n1213), .C(n1212), .D(n42), .Z(n930) );
  COND2X1 U866 ( .A(n44), .B(n1214), .C(n1213), .D(n42), .Z(n931) );
  COND2X1 U867 ( .A(n44), .B(n1215), .C(n1214), .D(n42), .Z(n932) );
  COND2X1 U868 ( .A(n44), .B(n1216), .C(n1215), .D(n42), .Z(n933) );
  COND2X1 U869 ( .A(n44), .B(n1217), .C(n1216), .D(n42), .Z(n934) );
  COND2X1 U870 ( .A(n44), .B(n1218), .C(n1217), .D(n42), .Z(n935) );
  COND2X1 U871 ( .A(n44), .B(n1219), .C(n1218), .D(n42), .Z(n936) );
  COND2X1 U872 ( .A(n44), .B(n1220), .C(n1219), .D(n42), .Z(n937) );
  COND2X1 U873 ( .A(n44), .B(n1221), .C(n1220), .D(n42), .Z(n938) );
  COND2X1 U874 ( .A(n44), .B(n1222), .C(n1221), .D(n42), .Z(n939) );
  COND2X1 U875 ( .A(n44), .B(n1223), .C(n1222), .D(n42), .Z(n940) );
  COND2X1 U876 ( .A(n44), .B(n1224), .C(n1223), .D(n42), .Z(n941) );
  COND2X1 U877 ( .A(n44), .B(n1225), .C(n1224), .D(n42), .Z(n942) );
  COND2X1 U878 ( .A(n44), .B(n1226), .C(n1225), .D(n42), .Z(n943) );
  COND2X1 U879 ( .A(n44), .B(n1227), .C(n1226), .D(n42), .Z(n944) );
  COND2X1 U880 ( .A(n44), .B(n1228), .C(n1227), .D(n42), .Z(n945) );
  CND2IX1 U906 ( .B(n1748), .A(n1731), .Z(n1229) );
  COND2X1 U907 ( .A(n36), .B(n1728), .C(n1256), .D(n33), .Z(n787) );
  COND2X1 U908 ( .A(n36), .B(n1231), .C(n1230), .D(n33), .Z(n947) );
  COND2X1 U909 ( .A(n36), .B(n1232), .C(n1231), .D(n33), .Z(n948) );
  COND2X1 U910 ( .A(n36), .B(n1233), .C(n1232), .D(n33), .Z(n949) );
  COND2X1 U911 ( .A(n36), .B(n1234), .C(n1233), .D(n33), .Z(n950) );
  COND2X1 U912 ( .A(n36), .B(n1235), .C(n1234), .D(n33), .Z(n951) );
  COND2X1 U913 ( .A(n36), .B(n1236), .C(n1235), .D(n33), .Z(n952) );
  COND2X1 U914 ( .A(n36), .B(n1237), .C(n1236), .D(n33), .Z(n953) );
  COND2X1 U915 ( .A(n36), .B(n1238), .C(n1237), .D(n33), .Z(n954) );
  COND2X1 U916 ( .A(n36), .B(n1239), .C(n1238), .D(n33), .Z(n955) );
  COND2X1 U917 ( .A(n36), .B(n1240), .C(n1239), .D(n33), .Z(n956) );
  COND2X1 U918 ( .A(n36), .B(n1241), .C(n1240), .D(n33), .Z(n957) );
  COND2X1 U919 ( .A(n36), .B(n1242), .C(n1241), .D(n33), .Z(n958) );
  COND2X1 U920 ( .A(n36), .B(n1243), .C(n1242), .D(n33), .Z(n959) );
  COND2X1 U921 ( .A(n36), .B(n1244), .C(n1243), .D(n33), .Z(n960) );
  COND2X1 U922 ( .A(n36), .B(n1245), .C(n1244), .D(n33), .Z(n961) );
  COND2X1 U923 ( .A(n36), .B(n1246), .C(n1245), .D(n33), .Z(n962) );
  COND2X1 U924 ( .A(n36), .B(n1247), .C(n1246), .D(n33), .Z(n963) );
  COND2X1 U925 ( .A(n36), .B(n1248), .C(n1247), .D(n33), .Z(n964) );
  COND2X1 U926 ( .A(n36), .B(n1249), .C(n1248), .D(n33), .Z(n965) );
  COND2X1 U927 ( .A(n36), .B(n1250), .C(n1249), .D(n33), .Z(n966) );
  COND2X1 U928 ( .A(n36), .B(n1251), .C(n1250), .D(n33), .Z(n967) );
  COND2X1 U929 ( .A(n36), .B(n1252), .C(n1251), .D(n33), .Z(n968) );
  COND2X1 U930 ( .A(n36), .B(n1253), .C(n1252), .D(n33), .Z(n969) );
  COND2X1 U932 ( .A(n36), .B(n1255), .C(n1254), .D(n33), .Z(n971) );
  CND2IX1 U960 ( .B(n1748), .A(n1722), .Z(n1256) );
  COND2X1 U961 ( .A(n27), .B(n1721), .C(n1285), .D(n24), .Z(n788) );
  COND2X1 U978 ( .A(n27), .B(n1274), .C(n24), .D(n1273), .Z(n989) );
  CND2IX1 U1018 ( .B(n1748), .A(n1714), .Z(n1285) );
  COND2X1 U1019 ( .A(n18), .B(n1713), .C(n1316), .D(n15), .Z(n789) );
  COND2X1 U1020 ( .A(n18), .B(n1287), .C(n15), .D(n1286), .Z(n1001) );
  COND2X1 U1021 ( .A(n18), .B(n1288), .C(n15), .D(n1287), .Z(n1002) );
  COND2X1 U1022 ( .A(n18), .B(n1289), .C(n15), .D(n1288), .Z(n1003) );
  COND2X1 U1023 ( .A(n18), .B(n1290), .C(n15), .D(n1289), .Z(n1004) );
  COND2X1 U1024 ( .A(n18), .B(n1291), .C(n15), .D(n1290), .Z(n1005) );
  COND2X1 U1025 ( .A(n18), .B(n1292), .C(n15), .D(n1291), .Z(n1006) );
  COND2X1 U1026 ( .A(n18), .B(n1293), .C(n15), .D(n1292), .Z(n1007) );
  COND2X1 U1027 ( .A(n18), .B(n1294), .C(n15), .D(n1293), .Z(n1008) );
  COND2X1 U1028 ( .A(n18), .B(n1295), .C(n15), .D(n1294), .Z(n1009) );
  COND2X1 U1029 ( .A(n18), .B(n1296), .C(n15), .D(n1295), .Z(n1010) );
  COND2X1 U1030 ( .A(n18), .B(n1297), .C(n15), .D(n1296), .Z(n1011) );
  COND2X1 U1031 ( .A(n18), .B(n1298), .C(n15), .D(n1297), .Z(n1012) );
  COND2X1 U1032 ( .A(n18), .B(n1299), .C(n15), .D(n1298), .Z(n1013) );
  COND2X1 U1033 ( .A(n18), .B(n1300), .C(n15), .D(n1299), .Z(n1014) );
  COND2X1 U1034 ( .A(n18), .B(n1301), .C(n15), .D(n1300), .Z(n1015) );
  COND2X1 U1035 ( .A(n18), .B(n1302), .C(n15), .D(n1301), .Z(n1016) );
  COND2X1 U1036 ( .A(n18), .B(n1303), .C(n15), .D(n1302), .Z(n1017) );
  COND2X1 U1037 ( .A(n18), .B(n1304), .C(n15), .D(n1303), .Z(n1018) );
  COND2X1 U1038 ( .A(n18), .B(n1305), .C(n15), .D(n1304), .Z(n1019) );
  COND2X1 U1039 ( .A(n18), .B(n1306), .C(n15), .D(n1305), .Z(n1020) );
  COND2X1 U1040 ( .A(n18), .B(n1307), .C(n15), .D(n1306), .Z(n1021) );
  COND2X1 U1041 ( .A(n18), .B(n1308), .C(n15), .D(n1307), .Z(n1022) );
  COND2X1 U1042 ( .A(n18), .B(n1309), .C(n15), .D(n1308), .Z(n1023) );
  COND2X1 U1043 ( .A(n18), .B(n1310), .C(n15), .D(n1309), .Z(n1024) );
  COND2X1 U1044 ( .A(n18), .B(n1311), .C(n15), .D(n1310), .Z(n1025) );
  COND2X1 U1045 ( .A(n18), .B(n1312), .C(n15), .D(n1311), .Z(n1026) );
  COND2X1 U1046 ( .A(n18), .B(n1313), .C(n15), .D(n1312), .Z(n1027) );
  COND2X1 U1047 ( .A(n18), .B(n1314), .C(n15), .D(n1313), .Z(n1028) );
  COND2X1 U1048 ( .A(n18), .B(n1315), .C(n15), .D(n1314), .Z(n1029) );
  CND2IX1 U1080 ( .B(n1748), .A(n1706), .Z(n1316) );
  CFD1QXL clk_r_REG0_S1 ( .D(n343), .CP(n1683), .Q(n1677) );
  CFD1QXL clk_r_REG11_S1 ( .D(n345), .CP(n1683), .Q(n1676) );
  CFD1QXL clk_r_REG6_S1 ( .D(n369), .CP(n1683), .Q(n1671) );
  CFD1QXL clk_r_REG10_S1 ( .D(n372), .CP(n1683), .Q(n1669) );
  CFD1QXL clk_r_REG52_S1 ( .D(n450), .CP(n1683), .Q(n1651) );
  CFD1QXL clk_r_REG30_S1 ( .D(n475), .CP(n1683), .Q(n1643) );
  CFD1QXL clk_r_REG12_S1 ( .D(n423), .CP(n1683), .Q(n1657) );
  CFD1QXL clk_r_REG13_S1 ( .D(n424), .CP(n1683), .Q(n1656) );
  CFD1QXL clk_r_REG27_S1 ( .D(n496), .CP(n1683), .Q(n1640) );
  CFD1QXL clk_r_REG45_S1 ( .D(n520), .CP(n1683), .Q(n1634) );
  CFD1QXL clk_r_REG88_S1 ( .D(n680), .CP(n1683), .Q(n1587) );
  CFD1QXL clk_r_REG92_S1 ( .D(n694), .CP(n1683), .Q(n1584) );
  CFD1QXL clk_r_REG76_S1 ( .D(n635), .CP(n1683), .Q(n1602) );
  CFD1QXL clk_r_REG74_S1 ( .D(n651), .CP(n1683), .Q(n1596) );
  CFD1QXL clk_r_REG96_S1 ( .D(n718), .CP(n1683), .Q(n1578) );
  CFD1QXL clk_r_REG94_S1 ( .D(n706), .CP(n1683), .Q(n1581) );
  CFD1QXL clk_r_REG85_S1 ( .D(n666), .CP(n1683), .Q(n1592) );
  CFD1QXL clk_r_REG102_S1 ( .D(n728), .CP(n1683), .Q(n1575) );
  CFD1QXL clk_r_REG104_S1 ( .D(n738), .CP(n1683), .Q(n1572) );
  CFD1QXL clk_r_REG3_S1 ( .D(n348), .CP(n1683), .Q(n1675) );
  CFD1QXL clk_r_REG113_S1 ( .D(n284), .CP(n1683), .Q(n1680) );
  CFD1QXL clk_r_REG111_S1 ( .D(n1546), .CP(n1683), .Q(n1682) );
  CFD1QXL clk_r_REG112_S1 ( .D(n285), .CP(n1683), .Q(n1679) );
  CFD1QXL clk_r_REG7_S1 ( .D(n370), .CP(n1683), .Q(n1670) );
  CFD1QXL clk_r_REG8_S1 ( .D(n395), .CP(n1683), .Q(n1666) );
  CFD1QXL clk_r_REG38_S1 ( .D(n447), .CP(n1683), .Q(n1653) );
  CFD1QXL clk_r_REG25_S1 ( .D(n474), .CP(n1683), .Q(n1644) );
  CFD1QXL clk_r_REG24_S1 ( .D(n473), .CP(n1683), .Q(n1645) );
  CFD1QXL clk_r_REG100_S1 ( .D(n454), .CP(n1683), .Q(n1649) );
  CFD1QXL clk_r_REG36_S1 ( .D(n421), .CP(n1683), .Q(n1659) );
  CFD1QXL clk_r_REG19_S1 ( .D(n425), .CP(n1683), .Q(n1655) );
  CFD1QXL clk_r_REG29_S1 ( .D(n498), .CP(n1683), .Q(n1638) );
  CFD1QXL clk_r_REG33_S1 ( .D(n522), .CP(n1683), .Q(n1632) );
  CFD1QXL clk_r_REG91_S1 ( .D(n693), .CP(n1683), .Q(n1585) );
  CFD1QXL clk_r_REG93_S1 ( .D(n705), .CP(n1683), .Q(n1582) );
  CFD1QXL clk_r_REG64_S1 ( .D(n620), .CP(n1683), .Q(n1606) );
  CFD1QXL clk_r_REG98_S1 ( .D(n720), .CP(n1683), .Q(n1577) );
  CFD1QXL clk_r_REG95_S1 ( .D(n717), .CP(n1683), .Q(n1579) );
  CFD1QXL clk_r_REG87_S1 ( .D(n679), .CP(n1683), .Q(n1588) );
  CFD1QXL clk_r_REG43_S1 ( .D(n540), .CP(n1683), .Q(n1627) );
  CFD1QXL clk_r_REG103_S1 ( .D(n737), .CP(n1683), .Q(n1573) );
  CFD1QXL clk_r_REG71_S1 ( .D(n582), .CP(n1683), .Q(n1616) );
  CFD1QXL clk_r_REG55_S1 ( .D(n562), .CP(n1683), .Q(n1621) );
  CFD1QXL clk_r_REG58_S1 ( .D(n602), .CP(n1683), .Q(n1611) );
  CFD1QXL clk_r_REG84_S1 ( .D(n665), .CP(n1683), .Q(n1593) );
  CFD1QXL clk_r_REG105_S1 ( .D(n745), .CP(n1683), .Q(n1568) );
  CFD1QXL clk_r_REG4_S1 ( .D(n393), .CP(n1683), .Q(n1668) );
  CFD1QXL clk_r_REG14_S1 ( .D(n397), .CP(n1683), .Q(n1664) );
  CFD1QXL clk_r_REG23_S1 ( .D(n420), .CP(n1683), .Q(n1660) );
  CFD1QXL clk_r_REG20_S1 ( .D(n426), .CP(n1683), .Q(n1654) );
  CFD1QXL clk_r_REG26_S1 ( .D(n495), .CP(n1683), .Q(n1641) );
  CFD1QXL clk_r_REG21_S1 ( .D(n452), .CP(n1683), .Q(n1650) );
  CFD1QXL clk_r_REG18_S1 ( .D(n458), .CP(n1683), .Q(n1648) );
  CFD1QXL clk_r_REG15_S1 ( .D(n398), .CP(n1683), .Q(n1663) );
  CFD1QXL clk_r_REG16_S1 ( .D(n400), .CP(n1683), .Q(n1662) );
  CFD1QXL clk_r_REG77_S1 ( .D(n636), .CP(n1683), .Q(n1601) );
  CFD1QXL clk_r_REG83_S1 ( .D(n682), .CP(n1683), .Q(n1586) );
  CFD1QXL clk_r_REG59_S1 ( .D(n541), .CP(n1683), .Q(n1626) );
  CFD1QXL clk_r_REG89_S1 ( .D(n696), .CP(n1683), .Q(n1583) );
  CFD1QXL clk_r_REG42_S1 ( .D(n539), .CP(n1683), .Q(n1628) );
  CFD1QXL clk_r_REG68_S1 ( .D(n622), .CP(n1683), .Q(n1604) );
  CFD1QXL clk_r_REG101_S1 ( .D(n727), .CP(n1683), .Q(n1576) );
  CFD1QXL clk_r_REG90_S1 ( .D(n708), .CP(n1683), .Q(n1580) );
  CFD1QXL clk_r_REG81_S1 ( .D(n668), .CP(n1683), .Q(n1590) );
  CFD1QXL clk_r_REG97_S1 ( .D(n730), .CP(n1683), .Q(n1574) );
  CFD1QXL clk_r_REG60_S1 ( .D(n542), .CP(n1683), .Q(n1625) );
  CFD1QXL clk_r_REG62_S1 ( .D(n584), .CP(n1683), .Q(n1614) );
  CFD1QXL clk_r_REG49_S1 ( .D(n564), .CP(n1683), .Q(n1619) );
  CFD1QXL clk_r_REG66_S1 ( .D(n604), .CP(n1683), .Q(n1609) );
  CFD1QXL clk_r_REG75_S1 ( .D(n652), .CP(n1683), .Q(n1595) );
  CFD1QXL clk_r_REG110_S1 ( .D(n282), .CP(n1683), .Q(n1681) );
  CFD1QXL clk_r_REG107_S1 ( .D(n744), .CP(n1683), .Q(n1569) );
  CFD1QXL clk_r_REG106_S1 ( .D(n743), .CP(n1683), .Q(n1570) );
  CFD1QXL clk_r_REG115_S1 ( .D(n286), .CP(n1683), .Q(n1678) );
  CFD1QX1 clk_r_REG48_S1 ( .D(n563), .CP(n1683), .Q(n1620) );
  CFD1QX1 clk_r_REG47_S1 ( .D(n524), .CP(n1683), .Q(n1630) );
  CFD1QX1 clk_r_REG69_S1 ( .D(n606), .CP(n1683), .Q(n1608) );
  CFD1QX1 clk_r_REG67_S1 ( .D(n621), .CP(n1683), .Q(n1605) );
  CFD1QX1 clk_r_REG78_S1 ( .D(n639), .CP(n1683), .Q(n1598) );
  CFD1QX1 clk_r_REG72_S1 ( .D(n637), .CP(n1683), .Q(n1600) );
  CFD1QX1 clk_r_REG54_S1 ( .D(n561), .CP(n1683), .Q(n1622) );
  CFD1QX2 clk_r_REG51_S1 ( .D(n544), .CP(n1683), .Q(n1623) );
  CFD1QX1 clk_r_REG57_S1 ( .D(n601), .CP(n1683), .Q(n1612) );
  CFD1QX2 clk_r_REG53_S1 ( .D(n586), .CP(n1683), .Q(n1613) );
  CFD1QX2 clk_r_REG50_S1 ( .D(n543), .CP(n1683), .Q(n1624) );
  CFD1QX4 clk_r_REG99_S1 ( .D(n526), .CP(n1683), .Q(n1629) );
  CFD1QX1 clk_r_REG28_S1 ( .D(n497), .CP(n1683), .Q(n1639) );
  CFD1QX2 clk_r_REG82_S1 ( .D(n654), .CP(n1683), .Q(n1594) );
  CFD1QX1 clk_r_REG63_S1 ( .D(n619), .CP(n1683), .Q(n1607) );
  CFD1QX1 clk_r_REG70_S1 ( .D(n581), .CP(n1683), .Q(n1617) );
  CFD1QX1 clk_r_REG80_S1 ( .D(n667), .CP(n1683), .Q(n1591) );
  CFD1QX1 clk_r_REG46_S1 ( .D(n523), .CP(n1683), .Q(n1631) );
  CFD1QX1 clk_r_REG32_S1 ( .D(n521), .CP(n1683), .Q(n1633) );
  CFD1QX1 clk_r_REG31_S1 ( .D(n476), .CP(n1683), .Q(n1642) );
  CFD1QX2 clk_r_REG34_S1 ( .D(n499), .CP(n1683), .Q(n1637) );
  CFD1QX1 clk_r_REG79_S1 ( .D(n640), .CP(n1683), .Q(n1597) );
  CFD1QXL clk_r_REG1_S1 ( .D(n367), .CP(n1683), .Q(n1673) );
  CFD1QXL clk_r_REG9_S1 ( .D(n396), .CP(n1683), .Q(n1665) );
  CFD1QXL clk_r_REG40_S1 ( .D(n471), .CP(n1683), .Q(n1647) );
  CFD1QXL clk_r_REG2_S1 ( .D(n368), .CP(n1683), .Q(n1672) );
  CFD1QXL clk_r_REG22_S1 ( .D(n419), .CP(n1683), .Q(n1661) );
  CFD1QXL clk_r_REG39_S1 ( .D(n448), .CP(n1683), .Q(n1652) );
  CFD1QXL clk_r_REG37_S1 ( .D(n422), .CP(n1683), .Q(n1658) );
  CFD1QXL clk_r_REG5_S1 ( .D(n394), .CP(n1683), .Q(n1667) );
  CFD1QXL clk_r_REG109_S1 ( .D(n751), .CP(n1683), .Q(n1567) );
  CFD1QXL clk_r_REG41_S1 ( .D(n472), .CP(n1683), .Q(n1646) );
  CFD1QXL clk_r_REG17_S1 ( .D(n366), .CP(n1683), .Q(n1674) );
  CFD1QX1 clk_r_REG117_S1 ( .D(n740), .CP(n1683), .Q(n1571) );
  CFD1QX2 clk_r_REG73_S1 ( .D(n638), .CP(n1683), .Q(n1599) );
  CFD1QX1 clk_r_REG35_S1 ( .D(n500), .CP(n1683), .Q(n1636) );
  CFD1QX2 clk_r_REG56_S1 ( .D(n566), .CP(n1683), .Q(n1618) );
  CFD1QX2 clk_r_REG108_S1 ( .D(n624), .CP(n1683), .Q(n1603) );
  CFD1QX1 clk_r_REG44_S1 ( .D(n519), .CP(n1683), .Q(n1635) );
  CFD1QX2 clk_r_REG65_S1 ( .D(n603), .CP(n1683), .Q(n1610) );
  CFD1QX2 clk_r_REG61_S1 ( .D(n583), .CP(n1683), .Q(n1615) );
  CFD1QX2 clk_r_REG86_S1 ( .D(n669), .CP(n1683), .Q(n1589) );
  CNR2X2 U1242 ( .A(n6), .B(n1317), .Z(n1031) );
  CNR2X2 U1243 ( .A(n6), .B(n1318), .Z(n1032) );
  CNR2X2 U1244 ( .A(n6), .B(n1319), .Z(n1033) );
  CNR2X2 U1245 ( .A(n6), .B(n1320), .Z(n1034) );
  CNR2X2 U1246 ( .A(n6), .B(n1321), .Z(n1035) );
  CNR2X2 U1247 ( .A(n6), .B(n1322), .Z(n1036) );
  CNR2X2 U1248 ( .A(n6), .B(n1323), .Z(n1037) );
  CNR2X2 U1249 ( .A(n6), .B(n1324), .Z(n1038) );
  CNR2X2 U1250 ( .A(n6), .B(n1325), .Z(n1039) );
  CNR2X2 U1251 ( .A(n6), .B(n1337), .Z(n1051) );
  CNR2X2 U1252 ( .A(n6), .B(n1338), .Z(n1052) );
  CNR2X2 U1253 ( .A(n6), .B(n1339), .Z(n1053) );
  CNR2X2 U1254 ( .A(n6), .B(n1340), .Z(n1054) );
  CNR2X2 U1255 ( .A(n6), .B(n1341), .Z(n1055) );
  CNR2X2 U1256 ( .A(n6), .B(n1342), .Z(n1056) );
  CNR2X2 U1257 ( .A(n6), .B(n1343), .Z(n1057) );
  CNR2X2 U1258 ( .A(n6), .B(n1344), .Z(n1058) );
  CNR2X2 U1259 ( .A(n6), .B(n1345), .Z(n1059) );
  CNR2X2 U1260 ( .A(n6), .B(n1346), .Z(n1060) );
  CNR2X2 U1261 ( .A(n6), .B(n1347), .Z(n1061) );
  CNR2X2 U1262 ( .A(n6), .B(n1336), .Z(n1050) );
  CNR2X2 U1263 ( .A(n6), .B(n1335), .Z(n1049) );
  CNR2X2 U1264 ( .A(n6), .B(n1334), .Z(n1048) );
  CNR2X2 U1265 ( .A(n6), .B(n1333), .Z(n1047) );
  CNR2X2 U1266 ( .A(n6), .B(n1332), .Z(n1046) );
  CNR2X2 U1267 ( .A(n6), .B(n1331), .Z(n1045) );
  CNR2X2 U1268 ( .A(n6), .B(n1330), .Z(n1044) );
  CNR2X2 U1269 ( .A(n6), .B(n1329), .Z(n1043) );
  CNR2X2 U1270 ( .A(n6), .B(n1328), .Z(n1042) );
  CNR2X2 U1271 ( .A(n6), .B(n1327), .Z(n1041) );
  CNR2X2 U1272 ( .A(n6), .B(n1326), .Z(n1040) );
  CIVX2 U1273 ( .A(b[28]), .Z(n1320) );
  CIVX2 U1274 ( .A(b[29]), .Z(n1319) );
  CIVX2 U1275 ( .A(b[27]), .Z(n1321) );
  CIVX2 U1276 ( .A(b[26]), .Z(n1322) );
  CIVX2 U1277 ( .A(b[24]), .Z(n1324) );
  CIVX2 U1278 ( .A(b[30]), .Z(n1318) );
  CIVX2 U1279 ( .A(b[25]), .Z(n1323) );
  CIVX2 U1280 ( .A(n1359), .Z(n1326) );
  CIVX2 U1281 ( .A(n1361), .Z(n1328) );
  CIVX2 U1282 ( .A(n1690), .Z(n1341) );
  CIVX2 U1283 ( .A(n1362), .Z(n1329) );
  CIVX2 U1284 ( .A(n1358), .Z(n1325) );
  CIVX2 U1285 ( .A(n1360), .Z(n1327) );
  CIVX2 U1286 ( .A(n1695), .Z(n1336) );
  CIVX2 U1287 ( .A(n1365), .Z(n1332) );
  CIVX2 U1288 ( .A(n1698), .Z(n1333) );
  CIVX2 U1289 ( .A(n1697), .Z(n1334) );
  CIVX2 U1290 ( .A(n1696), .Z(n1335) );
  CIVX2 U1291 ( .A(n1364), .Z(n1331) );
  CIVX2 U1292 ( .A(n1061), .Z(n308) );
  CIVX2 U1293 ( .A(n308), .Z(product[1]) );
  CIVX2 U1294 ( .A(n147), .Z(product[2]) );
  CIVX2 U1295 ( .A(n304), .Z(n302) );
  CIVX2 U1296 ( .A(a[2]), .Z(n15) );
  CIVX2 U1297 ( .A(b[31]), .Z(n1317) );
  CIVX2 U1298 ( .A(n1363), .Z(n1330) );
  CIVX2 U1299 ( .A(n1693), .Z(n1338) );
  CIVX2 U1300 ( .A(n1692), .Z(n1339) );
  CIVX2 U1301 ( .A(n1694), .Z(n1337) );
  CIVX2 U1302 ( .A(n1691), .Z(n1340) );
  CIVX2 U1303 ( .A(n1689), .Z(n1342) );
  CIVX2 U1304 ( .A(n1688), .Z(n1343) );
  CIVX2 U1305 ( .A(n1687), .Z(n1344) );
  CIVX2 U1306 ( .A(n1685), .Z(n1346) );
  CIVX2 U1307 ( .A(n1686), .Z(n1345) );
  CIVX2 U1308 ( .A(n1684), .Z(n1347) );
  CENXL U1309 ( .A(n1708), .B(n1686), .Z(n1312) );
  CND2XL U1310 ( .A(n1630), .B(n1624), .Z(n1527) );
  CND2XL U1311 ( .A(n1629), .B(n1630), .Z(n1525) );
  CANR1X1 U1312 ( .A(n257), .B(n265), .C(n258), .Z(n256) );
  CANR1X1 U1313 ( .A(n172), .B(n1552), .C(n167), .Z(n165) );
  CIVXL U1314 ( .A(n30), .Z(n1729) );
  CANR1XL U1315 ( .A(n201), .B(n1550), .C(n1522), .Z(n1519) );
  CANR1XL U1316 ( .A(n214), .B(n1551), .C(n209), .Z(n1520) );
  CIVX1 U1317 ( .A(n189), .Z(n187) );
  CANR1X1 U1318 ( .A(n214), .B(n1551), .C(n209), .Z(n207) );
  CND2XL U1319 ( .A(n1551), .B(n1558), .Z(n206) );
  CIVXL U1320 ( .A(n1522), .Z(n1521) );
  CAN2X1 U1321 ( .A(n556), .B(n575), .Z(n1522) );
  CND2X2 U1322 ( .A(n1533), .B(n1548), .Z(n179) );
  COND1X1 U1323 ( .A(n1534), .B(n1535), .C(n154), .Z(n1547) );
  CND2XL U1324 ( .A(n1550), .B(n1521), .Z(n127) );
  CANR1X1 U1325 ( .A(n201), .B(n1550), .C(n1522), .Z(n192) );
  CNR2X1 U1326 ( .A(n179), .B(n191), .Z(n177) );
  CEOX2 U1327 ( .A(n1709), .B(a[4]), .Z(n1564) );
  CENXL U1328 ( .A(n1709), .B(b[29]), .Z(n1286) );
  CENXL U1329 ( .A(n1709), .B(n1694), .Z(n1304) );
  CENXL U1330 ( .A(n1709), .B(n1684), .Z(n1314) );
  CIVX1 U1331 ( .A(n1713), .Z(n1709) );
  CIVX4 U1332 ( .A(n1564), .Z(n24) );
  CENX1 U1333 ( .A(n518), .B(n1523), .Z(n514) );
  CENX1 U1334 ( .A(n1628), .B(n537), .Z(n1523) );
  CIVXL U1335 ( .A(n221), .Z(n322) );
  COND1X2 U1336 ( .A(n278), .B(n266), .C(n267), .Z(n265) );
  CANR1X2 U1337 ( .A(n274), .B(n1563), .C(n269), .Z(n267) );
  CIVDX1 U1338 ( .A(n1749), .Z1(product[7]) );
  COND1X1 U1339 ( .A(n179), .B(n192), .C(n180), .Z(n178) );
  CENXL U1340 ( .A(n1692), .B(n1703), .Z(n1086) );
  CENXL U1341 ( .A(n1747), .B(n1703), .Z(n1095) );
  CENXL U1342 ( .A(n1688), .B(n1703), .Z(n1090) );
  CIVXL U1343 ( .A(n1703), .Z(n1411) );
  CENXL U1344 ( .A(n1687), .B(n1703), .Z(n1091) );
  CENXL U1345 ( .A(n1686), .B(n1703), .Z(n1092) );
  CENXL U1346 ( .A(n1684), .B(n1703), .Z(n1094) );
  CENXL U1347 ( .A(n1685), .B(n1703), .Z(n1093) );
  CENXL U1348 ( .A(n1689), .B(n1703), .Z(n1089) );
  CENXL U1349 ( .A(n1691), .B(n1703), .Z(n1087) );
  CENXL U1350 ( .A(n1690), .B(n1703), .Z(n1088) );
  CENX2 U1351 ( .A(n1703), .B(a[24]), .Z(n100) );
  CEO3X2 U1352 ( .A(n1629), .B(n1630), .C(n1624), .Z(n518) );
  CND2X1 U1353 ( .A(n1629), .B(n1624), .Z(n1526) );
  CND3X2 U1354 ( .A(n1525), .B(n1526), .C(n1527), .Z(n517) );
  CND2XL U1355 ( .A(n1628), .B(n537), .Z(n1528) );
  CND2XL U1356 ( .A(n1628), .B(n518), .Z(n1529) );
  CND2XL U1357 ( .A(n537), .B(n518), .Z(n1530) );
  CND3X1 U1358 ( .A(n1528), .B(n1529), .C(n1530), .Z(n513) );
  CIVX1 U1359 ( .A(n1713), .Z(n1712) );
  CIVX1 U1360 ( .A(n12), .Z(n1713) );
  COAN1X1 U1361 ( .A(n189), .B(n1531), .C(n184), .Z(n180) );
  CNR2XL U1362 ( .A(n512), .B(n533), .Z(n1531) );
  CIVDXL U1363 ( .A(n184), .Z0(n182) );
  COR2X2 U1364 ( .A(n512), .B(n533), .Z(n1533) );
  CIVXL U1365 ( .A(n182), .Z(n1532) );
  CNR2X1 U1366 ( .A(n384), .B(n411), .Z(n1534) );
  COAN1X1 U1367 ( .A(n156), .B(n158), .C(n157), .Z(n1535) );
  CND2XL U1368 ( .A(n384), .B(n411), .Z(n154) );
  COND1XL U1369 ( .A(n1519), .B(n179), .C(n180), .Z(n1536) );
  CENXL U1370 ( .A(n143), .B(n291), .Z(product[6]) );
  COND2XL U1371 ( .A(n27), .B(n1265), .C(n24), .D(n1264), .Z(n980) );
  COND2XL U1372 ( .A(n27), .B(n1279), .C(n24), .D(n1278), .Z(n994) );
  COND2XL U1373 ( .A(n27), .B(n1258), .C(n24), .D(n1257), .Z(n973) );
  COND2XL U1374 ( .A(n27), .B(n1260), .C(n24), .D(n1259), .Z(n975) );
  COND2XL U1375 ( .A(n27), .B(n1261), .C(n24), .D(n1260), .Z(n976) );
  COND2XL U1376 ( .A(n27), .B(n1262), .C(n24), .D(n1261), .Z(n977) );
  COND2XL U1377 ( .A(n27), .B(n1271), .C(n24), .D(n1270), .Z(n986) );
  COND2XL U1378 ( .A(n27), .B(n1267), .C(n24), .D(n1266), .Z(n982) );
  COND2XL U1379 ( .A(n27), .B(n1280), .C(n24), .D(n1279), .Z(n995) );
  COND2XL U1380 ( .A(n27), .B(n1270), .C(n24), .D(n1269), .Z(n985) );
  COND2XL U1381 ( .A(n27), .B(n1269), .C(n24), .D(n1268), .Z(n984) );
  COND2XL U1382 ( .A(n27), .B(n1264), .C(n24), .D(n1263), .Z(n979) );
  COND2XL U1383 ( .A(n27), .B(n1272), .C(n24), .D(n1271), .Z(n987) );
  COND2XL U1384 ( .A(n27), .B(n1266), .C(n24), .D(n1265), .Z(n981) );
  COND2XL U1385 ( .A(n27), .B(n1283), .C(n24), .D(n1282), .Z(n998) );
  COND2XL U1386 ( .A(n27), .B(n1282), .C(n24), .D(n1281), .Z(n997) );
  COND2XL U1387 ( .A(n27), .B(n1263), .C(n24), .D(n1262), .Z(n978) );
  COND2XL U1388 ( .A(n27), .B(n1278), .C(n24), .D(n1277), .Z(n993) );
  COND2XL U1389 ( .A(n27), .B(n1268), .C(n24), .D(n1267), .Z(n983) );
  COND2XL U1390 ( .A(n27), .B(n1284), .C(n24), .D(n1283), .Z(n999) );
  COND2XL U1391 ( .A(n27), .B(n1277), .C(n24), .D(n1276), .Z(n992) );
  COND2XL U1392 ( .A(n27), .B(n1273), .C(n24), .D(n1272), .Z(n988) );
  COND2XL U1393 ( .A(n27), .B(n1275), .C(n24), .D(n1274), .Z(n990) );
  COND2XL U1394 ( .A(n27), .B(n1276), .C(n24), .D(n1275), .Z(n991) );
  COND2XL U1395 ( .A(n27), .B(n1259), .C(n24), .D(n1258), .Z(n974) );
  COND2XL U1396 ( .A(n27), .B(n1281), .C(n24), .D(n1280), .Z(n996) );
  CIVX2 U1397 ( .A(n1730), .Z(n1727) );
  COND1X1 U1398 ( .A(n221), .B(n225), .C(n222), .Z(n220) );
  CANR1X2 U1399 ( .A(n234), .B(n1560), .C(n227), .Z(n225) );
  CENX4 U1400 ( .A(n1733), .B(a[10]), .Z(n50) );
  CIVX2 U1401 ( .A(n1739), .Z(n1733) );
  CANR1X1 U1402 ( .A(n238), .B(n219), .C(n220), .Z(n218) );
  CANR1XL U1403 ( .A(n205), .B(n177), .C(n1536), .Z(n1537) );
  COND1X1 U1404 ( .A(n206), .B(n218), .C(n207), .Z(n205) );
  COND1X1 U1405 ( .A(n256), .B(n239), .C(n240), .Z(n238) );
  COAN1XL U1406 ( .A(n206), .B(n218), .C(n1520), .Z(n1538) );
  CIVX1 U1407 ( .A(n1746), .Z(n1745) );
  CIVX2 U1408 ( .A(n55), .Z(n1746) );
  CEOX2 U1409 ( .A(n1718), .B(a[6]), .Z(n1561) );
  CENXL U1410 ( .A(n1718), .B(n1693), .Z(n1274) );
  CENXL U1411 ( .A(n1718), .B(n1691), .Z(n1276) );
  CENXL U1412 ( .A(n1718), .B(n1692), .Z(n1275) );
  CIVX3 U1413 ( .A(n1721), .Z(n1718) );
  CENXL U1414 ( .A(n149), .B(n1543), .Z(product[31]) );
  CIVXL U1415 ( .A(n163), .Z(n1539) );
  CIVX1 U1416 ( .A(n1539), .Z(n1540) );
  CENXL U1417 ( .A(n1540), .B(n122), .Z(product[27]) );
  CIVXL U1418 ( .A(n1537), .Z(n175) );
  CANR1X1 U1419 ( .A(n177), .B(n205), .C(n178), .Z(n176) );
  CANR1XL U1420 ( .A(n1553), .B(n1540), .C(n160), .Z(n1541) );
  COND1X1 U1421 ( .A(n164), .B(n176), .C(n165), .Z(n163) );
  COND2XL U1422 ( .A(n112), .B(n1067), .C(n110), .D(n1066), .Z(n794) );
  CNR2IXL U1423 ( .B(n1748), .A(n33), .Z(n972) );
  CND2X4 U1424 ( .A(n1391), .B(n58), .Z(n61) );
  CEOX1 U1425 ( .A(a[12]), .B(n1745), .Z(n1391) );
  CIVXL U1426 ( .A(n238), .Z(n237) );
  CNIVX1 U1427 ( .A(n1372), .Z(n1692) );
  CNR2X1 U1428 ( .A(n248), .B(n253), .Z(n246) );
  CNR2XL U1429 ( .A(n221), .B(n224), .Z(n219) );
  CIVX1 U1430 ( .A(n1743), .Z(n1742) );
  COND2X1 U1431 ( .A(n97), .B(n1089), .C(n1088), .D(n95), .Z(n813) );
  COR2XL U1432 ( .A(n1569), .B(n1567), .Z(n1562) );
  CAOR1XL U1433 ( .A(n238), .B(n219), .C(n220), .Z(n1542) );
  CANR1X1 U1434 ( .A(n1553), .B(n163), .C(n160), .Z(n158) );
  CNR2XL U1435 ( .A(n758), .B(n763), .Z(n284) );
  COND2XL U1436 ( .A(n69), .B(n1158), .C(n1157), .D(n66), .Z(n878) );
  COND2XL U1437 ( .A(n69), .B(n1156), .C(n1155), .D(n66), .Z(n876) );
  COND2X1 U1438 ( .A(n1076), .B(n105), .C(n1409), .D(n107), .Z(n777) );
  COND2X1 U1439 ( .A(n107), .B(n1073), .C(n105), .D(n1072), .Z(n799) );
  CND2X2 U1440 ( .A(n1390), .B(n66), .Z(n69) );
  CENX2 U1441 ( .A(n1741), .B(a[12]), .Z(n58) );
  CNIVX1 U1442 ( .A(n1379), .Z(n1685) );
  CND2IX4 U1443 ( .B(n1544), .A(n24), .Z(n27) );
  CNIVX1 U1444 ( .A(n1377), .Z(n1687) );
  CNIVX8 U1445 ( .A(n63), .Z(n1699) );
  CIVX2 U1446 ( .A(a[0]), .Z(n6) );
  CEOX1 U1447 ( .A(a[26]), .B(n1705), .Z(n1384) );
  CNIVX1 U1448 ( .A(n93), .Z(n1703) );
  CND2X1 U1449 ( .A(n95), .B(n1386), .Z(n97) );
  CNIVX4 U1450 ( .A(n86), .Z(n1702) );
  CND2X1 U1451 ( .A(n1385), .B(n100), .Z(n102) );
  CEOXL U1452 ( .A(n123), .B(n170), .Z(product[26]) );
  CND2XL U1453 ( .A(n1552), .B(n169), .Z(n123) );
  CND2XL U1454 ( .A(n312), .B(n157), .Z(n121) );
  CEOXL U1455 ( .A(n125), .B(n185), .Z(product[24]) );
  CND2XL U1456 ( .A(n1533), .B(n1532), .Z(n125) );
  CEOXL U1457 ( .A(n128), .B(n1538), .Z(product[21]) );
  CND2XL U1458 ( .A(n319), .B(n199), .Z(n128) );
  CND2XL U1459 ( .A(n1554), .B(n154), .Z(n120) );
  CND2XL U1460 ( .A(n1553), .B(n162), .Z(n122) );
  CND2XL U1461 ( .A(n1548), .B(n189), .Z(n126) );
  CND2XL U1462 ( .A(n1549), .B(n174), .Z(n124) );
  CND2XL U1463 ( .A(n319), .B(n1550), .Z(n191) );
  CND2XL U1464 ( .A(n752), .B(n757), .Z(n282) );
  CEOXL U1465 ( .A(n294), .B(n144), .Z(product[5]) );
  CNR2XL U1466 ( .A(n259), .B(n262), .Z(n257) );
  CND2XL U1467 ( .A(n1560), .B(n324), .Z(n224) );
  CEOXL U1468 ( .A(n129), .B(n212), .Z(product[20]) );
  CND2XL U1469 ( .A(n1551), .B(n211), .Z(n129) );
  CND2XL U1470 ( .A(n329), .B(n263), .Z(n138) );
  CND2XL U1471 ( .A(n1559), .B(n244), .Z(n134) );
  CND2XL U1472 ( .A(n324), .B(n232), .Z(n133) );
  CND2XL U1473 ( .A(n327), .B(n254), .Z(n136) );
  CND2XL U1474 ( .A(n1560), .B(n229), .Z(n132) );
  CND2XL U1475 ( .A(n322), .B(n222), .Z(n131) );
  CND2XL U1476 ( .A(n1558), .B(n216), .Z(n130) );
  COR2XL U1477 ( .A(n1060), .B(n1030), .Z(n1557) );
  COND2XL U1478 ( .A(n97), .B(n1088), .C(n1087), .D(n95), .Z(n812) );
  COND2XL U1479 ( .A(n84), .B(n1112), .C(n1111), .D(n82), .Z(n834) );
  COND2XL U1480 ( .A(n107), .B(n1071), .C(n105), .D(n1070), .Z(n797) );
  CNR2IXL U1481 ( .B(n1748), .A(n15), .Z(n1030) );
  CNR2IXL U1482 ( .B(n1748), .A(n74), .Z(n862) );
  CND2XL U1483 ( .A(n1563), .B(n271), .Z(n139) );
  CNR2IXL U1484 ( .B(n1748), .A(n114), .Z(n792) );
  CNR2IXL U1485 ( .B(n1748), .A(n82), .Z(n846) );
  CNR2IXL U1486 ( .B(n1748), .A(n95), .Z(n820) );
  COND2XL U1487 ( .A(n91), .B(n1107), .C(n1106), .D(n89), .Z(n830) );
  COND2XL U1488 ( .A(n102), .B(n1082), .C(n100), .D(n1081), .Z(n807) );
  CIVXL U1489 ( .A(n1705), .Z(n1409) );
  CNR2IXL U1490 ( .B(n1748), .A(n89), .Z(n832) );
  COND2XL U1491 ( .A(n84), .B(n1122), .C(n1121), .D(n82), .Z(n844) );
  CNR2IXL U1492 ( .B(n1748), .A(n105), .Z(n802) );
  COND2XL U1493 ( .A(n102), .B(n1083), .C(n100), .D(n1082), .Z(n808) );
  CNR2IXL U1494 ( .B(n1748), .A(n42), .Z(n946) );
  COND2XL U1495 ( .A(n36), .B(n1254), .C(n1253), .D(n33), .Z(n970) );
  CNR2IXL U1496 ( .B(n1748), .A(n100), .Z(n810) );
  COND2XL U1497 ( .A(n97), .B(n1094), .C(n1093), .D(n95), .Z(n818) );
  COND2XL U1498 ( .A(n112), .B(n1408), .C(n110), .D(n1069), .Z(n776) );
  COND2XL U1499 ( .A(n102), .B(n1080), .C(n100), .D(n1079), .Z(n805) );
  COND2XL U1500 ( .A(n84), .B(n1113), .C(n1112), .D(n82), .Z(n835) );
  CNR2IXL U1501 ( .B(n1748), .A(n110), .Z(n796) );
  COND2XL U1502 ( .A(n107), .B(n1074), .C(n105), .D(n1073), .Z(n800) );
  CND2XL U1503 ( .A(n716), .B(n725), .Z(n260) );
  CND2XL U1504 ( .A(n692), .B(n703), .Z(n249) );
  CND2IXL U1505 ( .B(n1748), .A(n1700), .Z(n1141) );
  CND2IXL U1506 ( .B(n1748), .A(n1703), .Z(n1096) );
  CND2IXL U1507 ( .B(n1748), .A(n1702), .Z(n1109) );
  CND2IXL U1508 ( .B(n1748), .A(n1704), .Z(n1085) );
  CND2IXL U1509 ( .B(n1748), .A(n1705), .Z(n1076) );
  CEOXL U1510 ( .A(n302), .B(n146), .Z(product[3]) );
  CND2XL U1511 ( .A(n1562), .B(n276), .Z(n140) );
  CNR2IXL U1512 ( .B(n1748), .A(n6), .Z(product[0]) );
  CENX1 U1513 ( .A(n340), .B(n355), .Z(n1543) );
  CENX2 U1514 ( .A(n1744), .B(a[14]), .Z(n66) );
  CENX2 U1515 ( .A(n1699), .B(a[16]), .Z(n74) );
  CNIVX2 U1516 ( .A(n99), .Z(n1704) );
  CNIVX4 U1517 ( .A(n71), .Z(n1700) );
  CND2X2 U1518 ( .A(n1388), .B(n82), .Z(n84) );
  CENXL U1519 ( .A(a[4]), .B(n1718), .Z(n1544) );
  CIVX3 U1520 ( .A(n1561), .Z(n33) );
  CND2IX2 U1521 ( .B(n1545), .A(n42), .Z(n44) );
  CENXL U1522 ( .A(a[8]), .B(n1737), .Z(n1545) );
  CNIVX1 U1523 ( .A(n1374), .Z(n1690) );
  CEOX1 U1524 ( .A(a[24]), .B(n1704), .Z(n1385) );
  CIVX3 U1525 ( .A(n1565), .Z(n42) );
  CND2XL U1526 ( .A(n1557), .B(n306), .Z(n147) );
  CND2IXL U1527 ( .B(n1748), .A(n113), .Z(n1064) );
  CND2IXL U1528 ( .B(n1748), .A(n109), .Z(n1069) );
  CIVXL U1529 ( .A(n109), .Z(n1408) );
  COND1XL U1530 ( .A(n191), .B(n1538), .C(n1519), .Z(n190) );
  CND2X1 U1531 ( .A(n1552), .B(n1549), .Z(n164) );
  COND1XL U1532 ( .A(n156), .B(n1541), .C(n157), .Z(n155) );
  COND1XL U1533 ( .A(n294), .B(n292), .C(n293), .Z(n291) );
  CENX1 U1534 ( .A(n197), .B(n127), .Z(product[22]) );
  COND1XL U1535 ( .A(n198), .B(n1538), .C(n199), .Z(n197) );
  CANR1XL U1536 ( .A(n291), .B(n1555), .C(n288), .Z(n286) );
  CND2X1 U1537 ( .A(n1555), .B(n290), .Z(n143) );
  CENX1 U1538 ( .A(n155), .B(n120), .Z(product[29]) );
  CENX1 U1539 ( .A(n190), .B(n126), .Z(product[23]) );
  CENX1 U1540 ( .A(n175), .B(n124), .Z(product[25]) );
  CND2X1 U1541 ( .A(n335), .B(n293), .Z(n144) );
  CEOXL U1542 ( .A(n121), .B(n1541), .Z(product[28]) );
  CANR1XL U1543 ( .A(n1549), .B(n175), .C(n172), .Z(n170) );
  CANR1XL U1544 ( .A(n1548), .B(n190), .C(n187), .Z(n185) );
  COR2X1 U1545 ( .A(n752), .B(n757), .Z(n1546) );
  CANR1XL U1546 ( .A(n299), .B(n1556), .C(n296), .Z(n294) );
  CANR1XL U1547 ( .A(n1558), .B(n1542), .C(n214), .Z(n212) );
  COND1XL U1548 ( .A(n263), .B(n259), .C(n260), .Z(n258) );
  CND2X1 U1549 ( .A(n246), .B(n1559), .Z(n239) );
  CANR1XL U1550 ( .A(n1559), .B(n247), .C(n242), .Z(n240) );
  COND1XL U1551 ( .A(n254), .B(n248), .C(n249), .Z(n247) );
  CENX1 U1552 ( .A(n145), .B(n299), .Z(product[4]) );
  CND2X1 U1553 ( .A(n1556), .B(n298), .Z(n145) );
  CENX1 U1554 ( .A(n261), .B(n137), .Z(product[12]) );
  CND2X1 U1555 ( .A(n328), .B(n260), .Z(n137) );
  COND1XL U1556 ( .A(n262), .B(n264), .C(n263), .Z(n261) );
  CENX1 U1557 ( .A(n255), .B(n136), .Z(product[13]) );
  CENX1 U1558 ( .A(n230), .B(n132), .Z(product[17]) );
  COND1XL U1559 ( .A(n231), .B(n237), .C(n232), .Z(n230) );
  CENX1 U1560 ( .A(n223), .B(n131), .Z(product[18]) );
  COND1XL U1561 ( .A(n224), .B(n237), .C(n225), .Z(n223) );
  CENX1 U1562 ( .A(n1542), .B(n130), .Z(product[19]) );
  CNR2X1 U1563 ( .A(n576), .B(n595), .Z(n198) );
  CNR2X1 U1564 ( .A(n412), .B(n437), .Z(n156) );
  CNR2X1 U1565 ( .A(n768), .B(n771), .Z(n292) );
  CNR2X1 U1566 ( .A(n774), .B(n789), .Z(n300) );
  CEOX1 U1567 ( .A(n138), .B(n264), .Z(product[11]) );
  CEOX1 U1568 ( .A(n135), .B(n250), .Z(product[14]) );
  CND2X1 U1569 ( .A(n326), .B(n249), .Z(n135) );
  CANR1XL U1570 ( .A(n327), .B(n255), .C(n252), .Z(n250) );
  CEOX1 U1571 ( .A(n134), .B(n245), .Z(product[15]) );
  CANR1XL U1572 ( .A(n246), .B(n255), .C(n247), .Z(n245) );
  CEOX1 U1573 ( .A(n133), .B(n237), .Z(product[16]) );
  COR2X1 U1574 ( .A(n534), .B(n555), .Z(n1548) );
  COR2X1 U1575 ( .A(n488), .B(n511), .Z(n1549) );
  COR2X1 U1576 ( .A(n575), .B(n556), .Z(n1550) );
  COR2X1 U1577 ( .A(n596), .B(n613), .Z(n1551) );
  CND2X1 U1578 ( .A(n576), .B(n595), .Z(n199) );
  COR2X1 U1579 ( .A(n464), .B(n487), .Z(n1552) );
  CND2X1 U1580 ( .A(n534), .B(n555), .Z(n189) );
  CND2X1 U1581 ( .A(n512), .B(n533), .Z(n184) );
  CND2X1 U1582 ( .A(n488), .B(n511), .Z(n174) );
  CND2X1 U1583 ( .A(n596), .B(n613), .Z(n211) );
  CND2X1 U1584 ( .A(n464), .B(n487), .Z(n169) );
  CND2X1 U1585 ( .A(n1060), .B(n1030), .Z(n306) );
  CND2X1 U1586 ( .A(n438), .B(n463), .Z(n162) );
  CND2X1 U1587 ( .A(n772), .B(n773), .Z(n298) );
  CND2X1 U1588 ( .A(n764), .B(n767), .Z(n290) );
  CND2X1 U1589 ( .A(n768), .B(n771), .Z(n293) );
  CND2XL U1590 ( .A(n774), .B(n789), .Z(n301) );
  CND2X1 U1591 ( .A(n412), .B(n437), .Z(n157) );
  COR2X1 U1592 ( .A(n438), .B(n463), .Z(n1553) );
  COR2X1 U1593 ( .A(n384), .B(n411), .Z(n1554) );
  COR2X1 U1594 ( .A(n764), .B(n767), .Z(n1555) );
  COR2X1 U1595 ( .A(n772), .B(n773), .Z(n1556) );
  CND2XL U1596 ( .A(n758), .B(n763), .Z(n285) );
  COND1XL U1597 ( .A(n302), .B(n300), .C(n301), .Z(n299) );
  CENX1 U1598 ( .A(n1702), .B(n1694), .Z(n1097) );
  CENX1 U1599 ( .A(n1700), .B(n1698), .Z(n1125) );
  CIVX2 U1600 ( .A(n1746), .Z(n1744) );
  CIVX2 U1601 ( .A(n1743), .Z(n1741) );
  CND2X1 U1602 ( .A(n1563), .B(n1562), .Z(n266) );
  CNR2X1 U1603 ( .A(n726), .B(n735), .Z(n262) );
  CNR2X1 U1604 ( .A(n632), .B(n647), .Z(n221) );
  CNR2X1 U1605 ( .A(n692), .B(n703), .Z(n248) );
  CNR2X1 U1606 ( .A(n716), .B(n725), .Z(n259) );
  CENX1 U1607 ( .A(n1733), .B(n1684), .Z(n1227) );
  CENX1 U1608 ( .A(n1741), .B(n1686), .Z(n1200) );
  CENX1 U1609 ( .A(n1744), .B(n1684), .Z(n1179) );
  CENX1 U1610 ( .A(n1744), .B(n1685), .Z(n1178) );
  CENX1 U1611 ( .A(n1699), .B(n1684), .Z(n1158) );
  CENX1 U1612 ( .A(n1744), .B(n1686), .Z(n1177) );
  CENX1 U1613 ( .A(n1734), .B(n1692), .Z(n1219) );
  CENX1 U1614 ( .A(n1725), .B(n1694), .Z(n1244) );
  CENX1 U1615 ( .A(n1736), .B(n1697), .Z(n1214) );
  CENX1 U1616 ( .A(n1702), .B(n1692), .Z(n1099) );
  CENX1 U1617 ( .A(n1723), .B(n1686), .Z(n1252) );
  CENX1 U1618 ( .A(n1723), .B(n1687), .Z(n1251) );
  CENX1 U1619 ( .A(n1733), .B(n1685), .Z(n1226) );
  CENX1 U1620 ( .A(n1725), .B(n1695), .Z(n1243) );
  CENX1 U1621 ( .A(n1735), .B(n1694), .Z(n1217) );
  CENX1 U1622 ( .A(n1726), .B(n1696), .Z(n1242) );
  CENX1 U1623 ( .A(n1734), .B(n1695), .Z(n1216) );
  CENX1 U1624 ( .A(n1735), .B(n1696), .Z(n1215) );
  CENX1 U1625 ( .A(n1736), .B(n1698), .Z(n1213) );
  CENX1 U1626 ( .A(n1725), .B(n1692), .Z(n1246) );
  CENX1 U1627 ( .A(n1724), .B(n1691), .Z(n1247) );
  CENX1 U1628 ( .A(n1723), .B(n1685), .Z(n1253) );
  CENX1 U1629 ( .A(n1724), .B(n1684), .Z(n1254) );
  CENX1 U1630 ( .A(n1732), .B(n1688), .Z(n1223) );
  CENX1 U1631 ( .A(n1732), .B(n1687), .Z(n1224) );
  CENX1 U1632 ( .A(n1732), .B(n1689), .Z(n1222) );
  CENX1 U1633 ( .A(n1734), .B(n1691), .Z(n1220) );
  CENX1 U1634 ( .A(n1732), .B(n1690), .Z(n1221) );
  CENX1 U1635 ( .A(n1725), .B(n1693), .Z(n1245) );
  CENX1 U1636 ( .A(n1726), .B(n1690), .Z(n1248) );
  CENX1 U1637 ( .A(n1722), .B(n1689), .Z(n1249) );
  CENX1 U1638 ( .A(n1723), .B(n1688), .Z(n1250) );
  CENX1 U1639 ( .A(n1726), .B(n1698), .Z(n1240) );
  CENX1 U1640 ( .A(n1733), .B(n1686), .Z(n1225) );
  CENX1 U1641 ( .A(n1726), .B(n1697), .Z(n1241) );
  CENX1 U1642 ( .A(n1741), .B(n1687), .Z(n1199) );
  CENX1 U1643 ( .A(n1741), .B(n1684), .Z(n1202) );
  CENX1 U1644 ( .A(n1741), .B(n1685), .Z(n1201) );
  CENX1 U1645 ( .A(n1741), .B(n1689), .Z(n1197) );
  CENX1 U1646 ( .A(n1741), .B(n1688), .Z(n1198) );
  CENX1 U1647 ( .A(n1699), .B(n1685), .Z(n1157) );
  CENX1 U1648 ( .A(n1744), .B(n1687), .Z(n1176) );
  CENX1 U1649 ( .A(n1741), .B(n1690), .Z(n1196) );
  CENX1 U1650 ( .A(n1699), .B(n1686), .Z(n1156) );
  CENX1 U1651 ( .A(n1700), .B(n1684), .Z(n1139) );
  CENX1 U1652 ( .A(n1744), .B(n1688), .Z(n1175) );
  CENX1 U1653 ( .A(n1699), .B(n1687), .Z(n1155) );
  CENX1 U1654 ( .A(n1741), .B(n1691), .Z(n1195) );
  CENX1 U1655 ( .A(n1744), .B(n1689), .Z(n1174) );
  CENX1 U1656 ( .A(n1700), .B(n1685), .Z(n1138) );
  CENX1 U1657 ( .A(n1701), .B(n1684), .Z(n1122) );
  CENX1 U1658 ( .A(n1700), .B(n1686), .Z(n1137) );
  CENX1 U1659 ( .A(n1744), .B(n1690), .Z(n1173) );
  CENX1 U1660 ( .A(n1699), .B(n1688), .Z(n1154) );
  CENX1 U1661 ( .A(n1744), .B(n1691), .Z(n1172) );
  CENX1 U1662 ( .A(n1700), .B(n1687), .Z(n1136) );
  CENX1 U1663 ( .A(n1699), .B(n1689), .Z(n1153) );
  CENX1 U1664 ( .A(n1701), .B(n1685), .Z(n1121) );
  CENX1 U1665 ( .A(n1744), .B(n1692), .Z(n1171) );
  CENX1 U1666 ( .A(n1700), .B(n1688), .Z(n1135) );
  CENX1 U1667 ( .A(n1699), .B(n1690), .Z(n1152) );
  CENX1 U1668 ( .A(n1684), .B(n1702), .Z(n1107) );
  CENX1 U1669 ( .A(n1702), .B(n1685), .Z(n1106) );
  CENX1 U1670 ( .A(n1701), .B(n1686), .Z(n1120) );
  CENX1 U1671 ( .A(n1742), .B(n1694), .Z(n1192) );
  CENX1 U1672 ( .A(n1699), .B(n1691), .Z(n1151) );
  CENX1 U1673 ( .A(n1701), .B(n1687), .Z(n1119) );
  CENX1 U1674 ( .A(n1742), .B(n1695), .Z(n1191) );
  CENX1 U1675 ( .A(n1744), .B(n1693), .Z(n1170) );
  CENX1 U1676 ( .A(n1700), .B(n1689), .Z(n1134) );
  CENX1 U1677 ( .A(n1699), .B(n1692), .Z(n1150) );
  CENX1 U1678 ( .A(n1701), .B(n1688), .Z(n1118) );
  CENX1 U1679 ( .A(n1702), .B(n1686), .Z(n1105) );
  CENX1 U1680 ( .A(n1702), .B(n1687), .Z(n1104) );
  CENX1 U1681 ( .A(n1744), .B(n1694), .Z(n1169) );
  CENX1 U1682 ( .A(n1700), .B(n1690), .Z(n1133) );
  CENX1 U1683 ( .A(n1744), .B(n1695), .Z(n1168) );
  CENX1 U1684 ( .A(n1700), .B(n1691), .Z(n1132) );
  CENX1 U1685 ( .A(n1699), .B(n1693), .Z(n1149) );
  CENX1 U1686 ( .A(n1701), .B(n1689), .Z(n1117) );
  CENX1 U1687 ( .A(n1699), .B(n1694), .Z(n1148) );
  CENX1 U1688 ( .A(n1701), .B(n1690), .Z(n1116) );
  CENX1 U1689 ( .A(n1742), .B(n1698), .Z(n1188) );
  CENX1 U1690 ( .A(n1700), .B(n1692), .Z(n1131) );
  CENX1 U1691 ( .A(n1702), .B(n1688), .Z(n1103) );
  CENX1 U1692 ( .A(n1745), .B(n1696), .Z(n1167) );
  CENX1 U1693 ( .A(n1699), .B(n1695), .Z(n1147) );
  CENX1 U1694 ( .A(n1702), .B(n1689), .Z(n1102) );
  CENX1 U1695 ( .A(n1745), .B(n1697), .Z(n1166) );
  CENX1 U1696 ( .A(n1700), .B(n1693), .Z(n1130) );
  CENX1 U1697 ( .A(n1700), .B(n1694), .Z(n1129) );
  CENX1 U1698 ( .A(n1699), .B(n1696), .Z(n1146) );
  CENX1 U1699 ( .A(n1702), .B(n1690), .Z(n1101) );
  CENX1 U1700 ( .A(n1745), .B(n1698), .Z(n1165) );
  CENX1 U1701 ( .A(n1701), .B(n1693), .Z(n1113) );
  CENX1 U1702 ( .A(n1700), .B(n1695), .Z(n1128) );
  CENX1 U1703 ( .A(n1702), .B(n1691), .Z(n1100) );
  CENX1 U1704 ( .A(n1699), .B(n1697), .Z(n1145) );
  CENX1 U1705 ( .A(n1700), .B(n1697), .Z(n1126) );
  CENX1 U1706 ( .A(n1700), .B(n1696), .Z(n1127) );
  CENX1 U1707 ( .A(n1702), .B(n1693), .Z(n1098) );
  CENX1 U1708 ( .A(n1699), .B(n1698), .Z(n1144) );
  CENX1 U1709 ( .A(n1701), .B(n1695), .Z(n1111) );
  CENX1 U1710 ( .A(n1701), .B(n1694), .Z(n1112) );
  CENX1 U1711 ( .A(n1735), .B(n1693), .Z(n1218) );
  CENX1 U1712 ( .A(n1742), .B(n1692), .Z(n1194) );
  CENX1 U1713 ( .A(n1742), .B(n1693), .Z(n1193) );
  CENX1 U1714 ( .A(n1741), .B(n1696), .Z(n1190) );
  CENX1 U1715 ( .A(n1742), .B(n1697), .Z(n1189) );
  CENX1 U1716 ( .A(n1701), .B(n1692), .Z(n1114) );
  CENX1 U1717 ( .A(n1701), .B(n1691), .Z(n1115) );
  CENX1 U1718 ( .A(n1717), .B(n1684), .Z(n1283) );
  CENX1 U1719 ( .A(n1710), .B(n1693), .Z(n1305) );
  CENX1 U1720 ( .A(n1710), .B(n1692), .Z(n1306) );
  CENX1 U1721 ( .A(n1711), .B(n1697), .Z(n1301) );
  CENX1 U1722 ( .A(n1711), .B(n1698), .Z(n1300) );
  CENX1 U1723 ( .A(n1719), .B(n1696), .Z(n1271) );
  CENX1 U1724 ( .A(n1719), .B(n1697), .Z(n1270) );
  CENX1 U1725 ( .A(n1720), .B(n1698), .Z(n1269) );
  CENX1 U1726 ( .A(n1717), .B(n1685), .Z(n1282) );
  CENX1 U1727 ( .A(n1716), .B(n1689), .Z(n1278) );
  CENX1 U1728 ( .A(n1716), .B(n1688), .Z(n1279) );
  CENX1 U1729 ( .A(n1710), .B(n1691), .Z(n1307) );
  CENX1 U1730 ( .A(n1708), .B(n1687), .Z(n1311) );
  CENX1 U1731 ( .A(n1708), .B(n1685), .Z(n1313) );
  CENX1 U1732 ( .A(n1711), .B(n1695), .Z(n1303) );
  CENX1 U1733 ( .A(n1711), .B(n1696), .Z(n1302) );
  CENX1 U1734 ( .A(n1708), .B(n1688), .Z(n1310) );
  CENX1 U1735 ( .A(n1719), .B(n1694), .Z(n1273) );
  CENX1 U1736 ( .A(n1707), .B(n1689), .Z(n1309) );
  CENX1 U1737 ( .A(n1707), .B(n1690), .Z(n1308) );
  CENX1 U1738 ( .A(n1717), .B(n1686), .Z(n1281) );
  CENX1 U1739 ( .A(n1716), .B(n1690), .Z(n1277) );
  CENX1 U1740 ( .A(n1716), .B(n1687), .Z(n1280) );
  CENX1 U1741 ( .A(n1719), .B(n1695), .Z(n1272) );
  CENX1 U1742 ( .A(n1684), .B(n1704), .Z(n1083) );
  CENX1 U1743 ( .A(n1685), .B(n1704), .Z(n1082) );
  CENX1 U1744 ( .A(n1686), .B(n1704), .Z(n1081) );
  CENX1 U1745 ( .A(n1687), .B(n1704), .Z(n1080) );
  CENX1 U1746 ( .A(n1685), .B(n1705), .Z(n1073) );
  CENX1 U1747 ( .A(n1686), .B(n1705), .Z(n1072) );
  CENX1 U1748 ( .A(n1689), .B(n1704), .Z(n1078) );
  CENX1 U1749 ( .A(n1688), .B(n1704), .Z(n1079) );
  CENX1 U1750 ( .A(n1687), .B(n1705), .Z(n1071) );
  CENX1 U1751 ( .A(n1684), .B(n1705), .Z(n1074) );
  CNR2X1 U1752 ( .A(n704), .B(n715), .Z(n253) );
  CENX1 U1753 ( .A(n1701), .B(n1696), .Z(n1110) );
  CENX1 U1754 ( .A(n1747), .B(n1727), .Z(n1255) );
  CENX1 U1755 ( .A(n1747), .B(n1737), .Z(n1228) );
  CENX1 U1756 ( .A(n1747), .B(n1742), .Z(n1203) );
  CENX1 U1757 ( .A(n1748), .B(n1745), .Z(n1180) );
  CENX1 U1758 ( .A(n1747), .B(n1699), .Z(n1159) );
  CENX1 U1759 ( .A(n1690), .B(n1704), .Z(n1077) );
  CENX1 U1760 ( .A(n1688), .B(n1705), .Z(n1070) );
  CENX1 U1761 ( .A(n1748), .B(n1700), .Z(n1140) );
  CENX1 U1762 ( .A(n1747), .B(n1701), .Z(n1123) );
  CENX1 U1763 ( .A(n1747), .B(n1702), .Z(n1108) );
  CENX1 U1764 ( .A(n1747), .B(n1704), .Z(n1084) );
  CENX1 U1765 ( .A(n1747), .B(n1705), .Z(n1075) );
  CNR2IX1 U1766 ( .B(n1748), .A(n24), .Z(n1000) );
  CENX1 U1767 ( .A(n1748), .B(n1720), .Z(n1284) );
  CENX1 U1768 ( .A(n1747), .B(n1712), .Z(n1315) );
  CNR2X1 U1769 ( .A(n664), .B(n677), .Z(n231) );
  CNR2IX1 U1770 ( .B(n1748), .A(n58), .Z(n900) );
  CND2XL U1771 ( .A(n337), .B(n301), .Z(n146) );
  COR2X1 U1772 ( .A(n614), .B(n631), .Z(n1558) );
  COR2X1 U1773 ( .A(n678), .B(n691), .Z(n1559) );
  COR2X1 U1774 ( .A(n648), .B(n663), .Z(n1560) );
  CND2X1 U1775 ( .A(n664), .B(n677), .Z(n232) );
  CND2X1 U1776 ( .A(n704), .B(n715), .Z(n254) );
  CNR2IX1 U1777 ( .B(n1748), .A(n66), .Z(n880) );
  CNR2IXL U1778 ( .B(n1748), .A(n50), .Z(n922) );
  CND2X1 U1779 ( .A(n726), .B(n735), .Z(n263) );
  CND2X1 U1780 ( .A(n648), .B(n663), .Z(n229) );
  CND2X1 U1781 ( .A(n614), .B(n631), .Z(n216) );
  CND2X1 U1782 ( .A(n678), .B(n691), .Z(n244) );
  CEOX1 U1783 ( .A(n797), .B(n811), .Z(n354) );
  CND2X1 U1784 ( .A(n632), .B(n647), .Z(n222) );
  CENX1 U1785 ( .A(n140), .B(n277), .Z(product[9]) );
  CEOX1 U1786 ( .A(n272), .B(n139), .Z(product[10]) );
  CANR1XL U1787 ( .A(n1562), .B(n277), .C(n274), .Z(n272) );
  CENX1 U1788 ( .A(n1704), .B(a[26]), .Z(n105) );
  CENX1 U1789 ( .A(n1700), .B(a[18]), .Z(n82) );
  CENX1 U1790 ( .A(n1701), .B(a[20]), .Z(n89) );
  CENX1 U1791 ( .A(n1705), .B(a[28]), .Z(n110) );
  CENX1 U1792 ( .A(n1702), .B(a[22]), .Z(n95) );
  COND1XL U1793 ( .A(n1680), .B(n1678), .C(n1679), .Z(n283) );
  CENX1 U1794 ( .A(n1734), .B(n1358), .Z(n1205) );
  CENX1 U1795 ( .A(n1724), .B(b[25]), .Z(n1230) );
  CENX1 U1796 ( .A(n109), .B(a[30]), .Z(n114) );
  CANR1XL U1797 ( .A(n1682), .B(n283), .C(n280), .Z(n278) );
  CEOX1 U1798 ( .A(a[2]), .B(n1712), .Z(n1396) );
  CEOX1 U1799 ( .A(a[6]), .B(n1727), .Z(n1394) );
  CENX1 U1800 ( .A(n1699), .B(n1364), .Z(n1142) );
  CENX1 U1801 ( .A(n1741), .B(n1360), .Z(n1182) );
  CENX1 U1802 ( .A(n1686), .B(n109), .Z(n1065) );
  CEOX1 U1803 ( .A(a[10]), .B(n1742), .Z(n1392) );
  CENX1 U1804 ( .A(n1741), .B(n1362), .Z(n1184) );
  CENX1 U1805 ( .A(n1745), .B(n1364), .Z(n1163) );
  CENX1 U1806 ( .A(n1742), .B(n1364), .Z(n1186) );
  CENX1 U1807 ( .A(n1736), .B(n1364), .Z(n1211) );
  CENX1 U1808 ( .A(n1722), .B(n1362), .Z(n1236) );
  CENX1 U1809 ( .A(n1727), .B(n1364), .Z(n1238) );
  CENX1 U1810 ( .A(n1731), .B(n1360), .Z(n1207) );
  CENX1 U1811 ( .A(n1726), .B(n1365), .Z(n1239) );
  CENX1 U1812 ( .A(n1727), .B(n1363), .Z(n1237) );
  CENX1 U1813 ( .A(n1731), .B(n1361), .Z(n1208) );
  CENX1 U1814 ( .A(n1736), .B(n1365), .Z(n1212) );
  CENX1 U1815 ( .A(n1735), .B(n1363), .Z(n1210) );
  CENX1 U1816 ( .A(n1722), .B(n1359), .Z(n1233) );
  CENX1 U1817 ( .A(n1731), .B(n1362), .Z(n1209) );
  CENX1 U1818 ( .A(n1722), .B(n1360), .Z(n1234) );
  CENX1 U1819 ( .A(n1731), .B(n1359), .Z(n1206) );
  CENX1 U1820 ( .A(n1726), .B(n1361), .Z(n1235) );
  CENX1 U1821 ( .A(n1722), .B(n1358), .Z(n1232) );
  CENX1 U1822 ( .A(n1745), .B(n1365), .Z(n1164) );
  CENX1 U1823 ( .A(n1742), .B(n1363), .Z(n1185) );
  CENX1 U1824 ( .A(n1745), .B(n1363), .Z(n1162) );
  CENX1 U1825 ( .A(n1699), .B(n1365), .Z(n1143) );
  CENX1 U1826 ( .A(n1741), .B(n1361), .Z(n1183) );
  CENX1 U1827 ( .A(n1722), .B(b[24]), .Z(n1231) );
  CENX1 U1828 ( .A(n1742), .B(n1365), .Z(n1187) );
  CENX1 U1829 ( .A(n1720), .B(n1364), .Z(n1267) );
  CENX1 U1830 ( .A(n1712), .B(n1364), .Z(n1298) );
  CENX1 U1831 ( .A(n1712), .B(n1365), .Z(n1299) );
  CENX1 U1832 ( .A(n1720), .B(n1365), .Z(n1268) );
  CENX1 U1833 ( .A(n1710), .B(n1363), .Z(n1297) );
  CENX1 U1834 ( .A(n1720), .B(n1363), .Z(n1266) );
  CENX1 U1835 ( .A(n1707), .B(n1361), .Z(n1295) );
  CENX1 U1836 ( .A(n1710), .B(n1359), .Z(n1293) );
  CENX1 U1837 ( .A(n1706), .B(n1358), .Z(n1292) );
  CENX1 U1838 ( .A(n1715), .B(n1359), .Z(n1262) );
  CENX1 U1839 ( .A(n1715), .B(n1358), .Z(n1261) );
  CENX1 U1840 ( .A(n1706), .B(b[26]), .Z(n1289) );
  CENX1 U1841 ( .A(n1714), .B(b[24]), .Z(n1260) );
  CENX1 U1842 ( .A(n1706), .B(b[27]), .Z(n1288) );
  CENX1 U1843 ( .A(n1706), .B(b[28]), .Z(n1287) );
  CENX1 U1844 ( .A(n1715), .B(n1361), .Z(n1264) );
  CENX1 U1845 ( .A(n1706), .B(b[25]), .Z(n1290) );
  CENX1 U1846 ( .A(n1710), .B(b[24]), .Z(n1291) );
  CENX1 U1847 ( .A(n1706), .B(n1362), .Z(n1296) );
  CENX1 U1848 ( .A(n1714), .B(n1362), .Z(n1265) );
  CENX1 U1849 ( .A(n1715), .B(n1360), .Z(n1263) );
  CENX1 U1850 ( .A(n1707), .B(n1360), .Z(n1294) );
  CENX1 U1851 ( .A(n1714), .B(b[25]), .Z(n1259) );
  CENX1 U1852 ( .A(n1714), .B(b[26]), .Z(n1258) );
  CENX1 U1853 ( .A(n1684), .B(n109), .Z(n1067) );
  CENX1 U1854 ( .A(n1685), .B(n109), .Z(n1066) );
  CEOXL U1855 ( .A(a[14]), .B(n1699), .Z(n1390) );
  CENX1 U1856 ( .A(n1745), .B(n1362), .Z(n1161) );
  CENX1 U1857 ( .A(n1717), .B(b[27]), .Z(n1257) );
  CENX1 U1858 ( .A(n1684), .B(n113), .Z(n1062) );
  CENX1 U1859 ( .A(n1747), .B(n113), .Z(n1063) );
  CENX1 U1860 ( .A(n1747), .B(n109), .Z(n1068) );
  CND2X2 U1861 ( .A(n1389), .B(n74), .Z(n77) );
  CEOXL U1862 ( .A(a[16]), .B(n1700), .Z(n1389) );
  CNIVX4 U1863 ( .A(n79), .Z(n1701) );
  CEOXL U1864 ( .A(a[18]), .B(n1701), .Z(n1388) );
  CNIVX1 U1865 ( .A(n116), .Z(n1747) );
  CNIVX2 U1866 ( .A(n1380), .Z(n1684) );
  CND2X1 U1867 ( .A(n89), .B(n1387), .Z(n91) );
  CEOXL U1868 ( .A(a[20]), .B(n1702), .Z(n1387) );
  CNIVX2 U1869 ( .A(n1378), .Z(n1686) );
  CND2X1 U1870 ( .A(n1384), .B(n105), .Z(n107) );
  CNIVX1 U1871 ( .A(n1376), .Z(n1688) );
  CNIVX1 U1872 ( .A(n1375), .Z(n1689) );
  COR2X1 U1873 ( .A(n736), .B(n1570), .Z(n1563) );
  CEOXL U1874 ( .A(a[22]), .B(n1703), .Z(n1386) );
  CNIVX1 U1875 ( .A(n116), .Z(n1748) );
  CNIVX1 U1876 ( .A(n1373), .Z(n1691) );
  CNIVX1 U1877 ( .A(n1371), .Z(n1693) );
  CNIVX1 U1878 ( .A(n1370), .Z(n1694) );
  CND2X1 U1879 ( .A(n736), .B(n1570), .Z(n271) );
  CND2X1 U1880 ( .A(n1569), .B(n1567), .Z(n276) );
  CND2X1 U1881 ( .A(n1383), .B(n110), .Z(n112) );
  CEOXL U1882 ( .A(a[28]), .B(n109), .Z(n1383) );
  CNIVX1 U1883 ( .A(n1369), .Z(n1695) );
  CNIVX1 U1884 ( .A(n1368), .Z(n1696) );
  CNIVX1 U1885 ( .A(n1367), .Z(n1697) );
  CNIVX1 U1886 ( .A(n1366), .Z(n1698) );
  CNIVX1 U1887 ( .A(n104), .Z(n1705) );
  CEOX1 U1888 ( .A(n1724), .B(a[8]), .Z(n1565) );
  CND2X1 U1889 ( .A(n1382), .B(n114), .Z(n115) );
  CEOXL U1890 ( .A(a[30]), .B(a[31]), .Z(n1382) );
  CENX1 U1891 ( .A(n141), .B(n283), .Z(product[8]) );
  CND2XL U1892 ( .A(n1682), .B(n1681), .Z(n141) );
  CEOXL U1893 ( .A(n1678), .B(n142), .Z(n1749) );
  CND2XL U1894 ( .A(n333), .B(n1679), .Z(n142) );
  CND2X4 U1895 ( .A(n1396), .B(n15), .Z(n18) );
  CND2X4 U1896 ( .A(n1394), .B(n33), .Z(n36) );
  CND2X4 U1897 ( .A(n1392), .B(n50), .Z(n53) );
  CIVXL U1898 ( .A(n1713), .Z(n1706) );
  CIVXL U1899 ( .A(n1713), .Z(n1707) );
  CIVXL U1900 ( .A(n1713), .Z(n1708) );
  CIVXL U1901 ( .A(n1713), .Z(n1710) );
  CIVXL U1902 ( .A(n1713), .Z(n1711) );
  CIVXL U1903 ( .A(n1721), .Z(n1714) );
  CIVXL U1904 ( .A(n1721), .Z(n1715) );
  CIVXL U1905 ( .A(n1721), .Z(n1716) );
  CIVXL U1906 ( .A(n1721), .Z(n1717) );
  CIVXL U1907 ( .A(n1721), .Z(n1719) );
  CIVXL U1908 ( .A(n1721), .Z(n1720) );
  CIVX2 U1909 ( .A(n21), .Z(n1721) );
  CIVXL U1910 ( .A(n1728), .Z(n1722) );
  CIVXL U1911 ( .A(n1729), .Z(n1723) );
  CIVXL U1912 ( .A(n1729), .Z(n1724) );
  CIVXL U1913 ( .A(n1730), .Z(n1725) );
  CIVXL U1914 ( .A(n1730), .Z(n1726) );
  CIVXL U1915 ( .A(n30), .Z(n1728) );
  CIVXL U1916 ( .A(n30), .Z(n1730) );
  CIVXL U1917 ( .A(n1738), .Z(n1731) );
  CIVXL U1918 ( .A(n1739), .Z(n1732) );
  CIVXL U1919 ( .A(n1739), .Z(n1734) );
  CIVXL U1920 ( .A(n1740), .Z(n1735) );
  CIVXL U1921 ( .A(n1740), .Z(n1736) );
  CIVXL U1922 ( .A(n1740), .Z(n1737) );
  CIVXL U1923 ( .A(n39), .Z(n1738) );
  CIVXL U1924 ( .A(n39), .Z(n1739) );
  CIVXL U1925 ( .A(n39), .Z(n1740) );
  CIVX1 U1926 ( .A(n48), .Z(n1743) );
  CIVX2 U1927 ( .A(n300), .Z(n337) );
  CIVX2 U1928 ( .A(n292), .Z(n335) );
  CIVX2 U1929 ( .A(n1680), .Z(n333) );
  CIVX2 U1930 ( .A(n262), .Z(n329) );
  CIVX2 U1931 ( .A(n259), .Z(n328) );
  CIVX2 U1932 ( .A(n248), .Z(n326) );
  CIVX2 U1933 ( .A(n156), .Z(n312) );
  CIVX2 U1934 ( .A(n306), .Z(n304) );
  CIVX2 U1935 ( .A(n298), .Z(n296) );
  CIVX2 U1936 ( .A(n290), .Z(n288) );
  CIVX2 U1937 ( .A(n1681), .Z(n280) );
  CIVX2 U1938 ( .A(n278), .Z(n277) );
  CIVX2 U1939 ( .A(n276), .Z(n274) );
  CIVX2 U1940 ( .A(n271), .Z(n269) );
  CIVX2 U1941 ( .A(n265), .Z(n264) );
  CIVX2 U1942 ( .A(n256), .Z(n255) );
  CIVX2 U1943 ( .A(n254), .Z(n252) );
  CIVX2 U1944 ( .A(n253), .Z(n327) );
  CIVX2 U1945 ( .A(n244), .Z(n242) );
  CIVX2 U1946 ( .A(n232), .Z(n234) );
  CIVX2 U1947 ( .A(n231), .Z(n324) );
  CIVX2 U1948 ( .A(n229), .Z(n227) );
  CIVX2 U1949 ( .A(n216), .Z(n214) );
  CIVX2 U1950 ( .A(n211), .Z(n209) );
  CIVX2 U1951 ( .A(n199), .Z(n201) );
  CIVX2 U1952 ( .A(n198), .Z(n319) );
  CIVX2 U1953 ( .A(n174), .Z(n172) );
  CIVX2 U1954 ( .A(n169), .Z(n167) );
  CIVX2 U1955 ( .A(n162), .Z(n160) );
  CIVX2 U1956 ( .A(n1699), .Z(n1415) );
  CIVX2 U1957 ( .A(n1700), .Z(n1414) );
  CIVX2 U1958 ( .A(n1701), .Z(n1413) );
  CIVX2 U1959 ( .A(n1702), .Z(n1412) );
  CIVX2 U1960 ( .A(n1704), .Z(n1410) );
  CIVX2 U1961 ( .A(n113), .Z(n1407) );
endmodule


module calc_DW02_mult_2_stage_3 ( A, B, TC, CLK, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC, CLK;
  wire   n27, n28, n29, n30, n31, n32, n33, \A_extended[32] , \B_extended[32] ,
         n7, n9, n11, n13, n15, n17, n19, n20, n21, n22, n23, n24, n25, n26;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33;
  assign \A_extended[32]  = A[31];
  assign \B_extended[32]  = B[31];

  calc_DW_mult_tc_18 mult_96 ( .a({\A_extended[32] , \A_extended[32] , A[30:2], 
        1'b0, A[0]}), .b({\B_extended[32] , \B_extended[32] , B[30:0]}), 
        .product({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, PRODUCT[31:7], n27, 
        n28, n29, n30, n31, n32, n33}), .dw8_CLK(CLK) );
  CFD1QXL clk_r_REG120_S1 ( .D(n31), .CP(CLK), .Q(n22) );
  CFD1QXL clk_r_REG121_S1 ( .D(n32), .CP(CLK), .Q(n21) );
  CFD1QXL clk_r_REG119_S1 ( .D(n30), .CP(CLK), .Q(n23) );
  CFD1QXL clk_r_REG122_S1 ( .D(n33), .CP(CLK), .Q(n20) );
  CFD1QXL clk_r_REG118_S1 ( .D(n29), .CP(CLK), .Q(n24) );
  CFD1QXL clk_r_REG114_S1 ( .D(n27), .CP(CLK), .Q(n26) );
  CFD1QXL clk_r_REG116_S1 ( .D(n28), .CP(CLK), .Q(n25) );
  CIVDXL U2 ( .A(n26), .Z1(n7) );
  CNIVX1 U3 ( .A(n7), .Z(PRODUCT[6]) );
  CIVDXL U4 ( .A(n22), .Z1(n9) );
  CNIVX1 U5 ( .A(n9), .Z(PRODUCT[2]) );
  CIVDXL U6 ( .A(n25), .Z1(n11) );
  CNIVX1 U7 ( .A(n11), .Z(PRODUCT[5]) );
  CIVDXL U8 ( .A(n24), .Z1(n13) );
  CNIVX1 U9 ( .A(n13), .Z(PRODUCT[4]) );
  CIVDXL U10 ( .A(n23), .Z1(n15) );
  CNIVX1 U11 ( .A(n15), .Z(PRODUCT[3]) );
  CIVDXL U12 ( .A(n20), .Z1(n17) );
  CNIVX1 U13 ( .A(n17), .Z(PRODUCT[0]) );
  CIVDXL U14 ( .A(n21), .Z1(n19) );
  CNIVX1 U15 ( .A(n19), .Z(PRODUCT[1]) );
endmodule


module calc_DW_mult_tc_16 ( a, b, product, dw6_CLK );
  input [32:0] a;
  input [32:0] b;
  output [65:0] product;
  input dw6_CLK;
  wire   n3, n6, n9, n12, n15, n18, n21, n24, n27, n30, n33, n36, n39, n42,
         n44, n48, n50, n53, n55, n58, n61, n63, n66, n69, n71, n74, n77, n79,
         n82, n84, n86, n89, n91, n93, n95, n97, n99, n100, n102, n104, n105,
         n107, n109, n110, n112, n113, n114, n115, n116, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n150, n151, n152, n153, n155, n157, n158,
         n159, n160, n161, n163, n165, n166, n167, n168, n170, n172, n173,
         n175, n177, n178, n179, n180, n181, n182, n183, n185, n187, n188,
         n190, n192, n193, n194, n195, n197, n199, n200, n201, n202, n204,
         n208, n209, n210, n212, n214, n215, n217, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n230, n232, n233, n234, n235,
         n237, n240, n241, n242, n243, n245, n247, n248, n249, n250, n251,
         n252, n253, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n272, n274, n275, n277,
         n279, n280, n281, n283, n285, n286, n287, n288, n289, n291, n293,
         n294, n295, n296, n297, n299, n301, n302, n303, n304, n305, n307,
         n309, n310, n312, n313, n315, n322, n325, n327, n329, n330, n331,
         n332, n336, n338, n340, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1395, n1396, n1397, n1399,
         n1400, n1410, n1411, n1412, n1766, n1765, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764;
  assign n3 = a[1];
  assign n12 = a[3];
  assign n21 = a[5];
  assign n30 = a[7];
  assign n39 = a[9];
  assign n48 = a[11];
  assign n55 = a[13];
  assign n63 = a[15];
  assign n71 = a[17];
  assign n79 = a[19];
  assign n86 = a[21];
  assign n93 = a[23];
  assign n99 = a[25];
  assign n104 = a[27];
  assign n109 = a[29];
  assign n113 = a[32];
  assign n116 = b[0];
  assign n1361 = b[23];
  assign n1362 = b[22];
  assign n1363 = b[21];
  assign n1364 = b[20];
  assign n1365 = b[19];
  assign n1366 = b[18];
  assign n1367 = b[17];
  assign n1368 = b[16];
  assign n1369 = b[15];
  assign n1370 = b[14];
  assign n1371 = b[13];
  assign n1372 = b[12];
  assign n1373 = b[11];
  assign n1374 = b[10];
  assign n1375 = b[9];
  assign n1376 = b[8];
  assign n1377 = b[7];
  assign n1378 = b[6];
  assign n1379 = b[5];
  assign n1380 = b[4];
  assign n1381 = b[3];
  assign n1382 = b[2];
  assign n1383 = b[1];
  assign n1692 = dw6_CLK;

  CEO3X2 U350 ( .A(n362), .B(n344), .C(n360), .Z(n343) );
  CEO3X2 U351 ( .A(n364), .B(n346), .C(n345), .Z(n344) );
  CEO3X2 U352 ( .A(n1684), .B(n366), .C(n347), .Z(n345) );
  CEO3X2 U353 ( .A(n1678), .B(n1680), .C(n1683), .Z(n346) );
  CEO3X2 U354 ( .A(n1676), .B(n1681), .C(n1682), .Z(n347) );
  CEO3X2 U355 ( .A(n353), .B(n352), .C(n374), .Z(n348) );
  CEO3X2 U356 ( .A(n356), .B(n355), .C(n354), .Z(n349) );
  CEO3X2 U357 ( .A(n380), .B(n376), .C(n378), .Z(n350) );
  CEO3X2 U358 ( .A(n357), .B(n384), .C(n382), .Z(n351) );
  CEO3X2 U359 ( .A(n926), .B(n950), .C(n1034), .Z(n352) );
  CEO3X2 U360 ( .A(n904), .B(n976), .C(n1004), .Z(n353) );
  CEO3X2 U361 ( .A(n794), .B(n866), .C(n884), .Z(n354) );
  CEO3X2 U362 ( .A(n814), .B(n824), .C(n850), .Z(n355) );
  CEO3X2 U363 ( .A(n800), .B(n796), .C(n836), .Z(n356) );
  CFA1X1 U365 ( .A(n363), .B(n361), .CI(n388), .CO(n358), .S(n359) );
  CFA1X1 U366 ( .A(n367), .B(n390), .CI(n365), .CO(n360), .S(n361) );
  CFA1X1 U367 ( .A(n1679), .B(n392), .CI(n394), .CO(n362), .S(n363) );
  CFA1X1 U368 ( .A(n1673), .B(n1677), .CI(n1675), .CO(n364), .S(n365) );
  CFA1X1 U369 ( .A(n1669), .B(n1674), .CI(n1671), .CO(n366), .S(n367) );
  CFA1X1 U370 ( .A(n402), .B(n377), .CI(n379), .CO(n368), .S(n369) );
  CFA1X1 U371 ( .A(n385), .B(n381), .CI(n383), .CO(n370), .S(n371) );
  CFA1X1 U372 ( .A(n410), .B(n404), .CI(n406), .CO(n372), .S(n373) );
  CFA1X1 U373 ( .A(n927), .B(n408), .CI(n412), .CO(n374), .S(n375) );
  CFA1X1 U374 ( .A(n905), .B(n1035), .CI(n951), .CO(n376), .S(n377) );
  CFA1X1 U375 ( .A(n885), .B(n977), .CI(n1005), .CO(n378), .S(n379) );
  CFA1X1 U376 ( .A(n797), .B(n867), .CI(n837), .CO(n380), .S(n381) );
  CFA1X1 U377 ( .A(n801), .B(n851), .CI(n825), .CO(n382), .S(n383) );
  CFA1X1 U378 ( .A(n795), .B(n815), .CI(n807), .CO(n384), .S(n385) );
  CFA1X1 U379 ( .A(n391), .B(n389), .CI(n416), .CO(n386), .S(n387) );
  CFA1X1 U380 ( .A(n395), .B(n418), .CI(n393), .CO(n388), .S(n389) );
  CFA1X1 U381 ( .A(n1672), .B(n420), .CI(n422), .CO(n390), .S(n391) );
  CFA1X1 U382 ( .A(n1668), .B(n1670), .CI(n1666), .CO(n392), .S(n393) );
  CFA1X1 U383 ( .A(n1667), .B(n1664), .CI(n1662), .CO(n394), .S(n395) );
  CFA1X1 U384 ( .A(n409), .B(n405), .CI(n407), .CO(n396), .S(n397) );
  CFA1X1 U385 ( .A(n430), .B(n411), .CI(n432), .CO(n398), .S(n399) );
  CFA1X1 U386 ( .A(n438), .B(n434), .CI(n436), .CO(n400), .S(n401) );
  CFA1X1 U387 ( .A(n928), .B(n413), .CI(n952), .CO(n402), .S(n403) );
  CFA1X1 U388 ( .A(n906), .B(n978), .CI(n1036), .CO(n404), .S(n405) );
  CFA1X1 U389 ( .A(n838), .B(n1006), .CI(n886), .CO(n406), .S(n407) );
  CFA1X1 U390 ( .A(n816), .B(n868), .CI(n798), .CO(n408), .S(n409) );
  CFA1X1 U391 ( .A(n802), .B(n852), .CI(n826), .CO(n410), .S(n411) );
  CHA1X1 U392 ( .A(n779), .B(n808), .CO(n412), .S(n413) );
  CFA1X1 U393 ( .A(n419), .B(n417), .CI(n442), .CO(n414), .S(n415) );
  CFA1X1 U394 ( .A(n423), .B(n444), .CI(n421), .CO(n416), .S(n417) );
  CFA1X1 U395 ( .A(n1665), .B(n446), .CI(n448), .CO(n418), .S(n419) );
  CFA1X1 U396 ( .A(n1661), .B(n1663), .CI(n1659), .CO(n420), .S(n421) );
  CFA1X1 U397 ( .A(n1660), .B(n1657), .CI(n1655), .CO(n422), .S(n423) );
  CFA1X1 U398 ( .A(n437), .B(n433), .CI(n435), .CO(n424), .S(n425) );
  CFA1X1 U399 ( .A(n458), .B(n439), .CI(n456), .CO(n426), .S(n427) );
  CFA1X1 U400 ( .A(n464), .B(n462), .CI(n460), .CO(n428), .S(n429) );
  CFA1X1 U401 ( .A(n907), .B(n953), .CI(n929), .CO(n430), .S(n431) );
  CFA1X1 U402 ( .A(n887), .B(n979), .CI(n1037), .CO(n432), .S(n433) );
  CFA1X1 U403 ( .A(n839), .B(n1007), .CI(n853), .CO(n434), .S(n435) );
  CFA1X1 U404 ( .A(n803), .B(n869), .CI(n827), .CO(n436), .S(n437) );
  CFA1X1 U405 ( .A(n799), .B(n817), .CI(n809), .CO(n438), .S(n439) );
  CFA1X1 U406 ( .A(n445), .B(n443), .CI(n468), .CO(n440), .S(n441) );
  CFA1X1 U407 ( .A(n449), .B(n470), .CI(n447), .CO(n442), .S(n443) );
  CFA1X1 U408 ( .A(n1651), .B(n472), .CI(n1658), .CO(n444), .S(n445) );
  CFA1X1 U409 ( .A(n1654), .B(n1656), .CI(n1649), .CO(n446), .S(n447) );
  CFA1X1 U410 ( .A(n1652), .B(n1647), .CI(n1653), .CO(n448), .S(n449) );
  CFA1X1 U411 ( .A(n480), .B(n459), .CI(n461), .CO(n450), .S(n451) );
  CFA1X1 U412 ( .A(n486), .B(n482), .CI(n484), .CO(n452), .S(n453) );
  CFA1X1 U413 ( .A(n954), .B(n488), .CI(n465), .CO(n454), .S(n455) );
  CFA1X1 U414 ( .A(n930), .B(n1008), .CI(n1038), .CO(n456), .S(n457) );
  CFA1X1 U415 ( .A(n854), .B(n980), .CI(n908), .CO(n458), .S(n459) );
  CFA1X1 U416 ( .A(n828), .B(n870), .CI(n818), .CO(n460), .S(n461) );
  CFA1X1 U417 ( .A(n804), .B(n888), .CI(n840), .CO(n462), .S(n463) );
  CHA1X1 U418 ( .A(n780), .B(n810), .CO(n464), .S(n465) );
  CFA1X1 U419 ( .A(n471), .B(n469), .CI(n492), .CO(n466), .S(n467) );
  CFA1X1 U420 ( .A(n496), .B(n494), .CI(n473), .CO(n468), .S(n469) );
  CFA1X1 U421 ( .A(n1645), .B(n1650), .CI(n1648), .CO(n470), .S(n471) );
  CFA1X1 U422 ( .A(n1641), .B(n1646), .CI(n1643), .CO(n472), .S(n473) );
  CFA1X1 U423 ( .A(n485), .B(n481), .CI(n483), .CO(n474), .S(n475) );
  CFA1X1 U424 ( .A(n506), .B(n487), .CI(n489), .CO(n476), .S(n477) );
  CFA1X1 U425 ( .A(n510), .B(n504), .CI(n508), .CO(n478), .S(n479) );
  CFA1X1 U426 ( .A(n931), .B(n512), .CI(n955), .CO(n480), .S(n481) );
  CFA1X1 U427 ( .A(n871), .B(n981), .CI(n1039), .CO(n482), .S(n483) );
  CFA1X1 U429 ( .A(n829), .B(n889), .CI(n841), .CO(n486), .S(n487) );
  CFA1X1 U430 ( .A(n805), .B(n811), .CI(n819), .CO(n488), .S(n489) );
  CFA1X1 U431 ( .A(n495), .B(n493), .CI(n516), .CO(n490), .S(n491) );
  CFA1X1 U432 ( .A(n520), .B(n518), .CI(n497), .CO(n492), .S(n493) );
  CFA1X1 U433 ( .A(n1639), .B(n1644), .CI(n1642), .CO(n494), .S(n495) );
  CFA1X1 U434 ( .A(n1635), .B(n1640), .CI(n1637), .CO(n496), .S(n497) );
  CFA1X1 U435 ( .A(n509), .B(n505), .CI(n507), .CO(n498), .S(n499) );
  CFA1X1 U436 ( .A(n530), .B(n511), .CI(n528), .CO(n500), .S(n501) );
  CFA1X1 U437 ( .A(n513), .B(n532), .CI(n534), .CO(n502), .S(n503) );
  CFA1X1 U438 ( .A(n932), .B(n1010), .CI(n956), .CO(n504), .S(n505) );
  CFA1X1 U439 ( .A(n872), .B(n982), .CI(n1040), .CO(n506), .S(n507) );
  CFA1X1 U441 ( .A(n820), .B(n910), .CI(n842), .CO(n510), .S(n511) );
  CHA1X1 U442 ( .A(n781), .B(n812), .CO(n512), .S(n513) );
  CFA1X1 U443 ( .A(n519), .B(n517), .CI(n538), .CO(n514), .S(n515) );
  CFA1X1 U444 ( .A(n542), .B(n521), .CI(n540), .CO(n516), .S(n517) );
  CFA1X1 U445 ( .A(n1632), .B(n1638), .CI(n1636), .CO(n518), .S(n519) );
  CFA1X1 U446 ( .A(n1633), .B(n1634), .CI(n1630), .CO(n520), .S(n521) );
  CFA1X1 U447 ( .A(n533), .B(n548), .CI(n531), .CO(n522), .S(n523) );
  CFA1X1 U448 ( .A(n554), .B(n535), .CI(n550), .CO(n524), .S(n525) );
  CFA1X1 U449 ( .A(n933), .B(n552), .CI(n556), .CO(n526), .S(n527) );
  CFA1X1 U450 ( .A(n891), .B(n1041), .CI(n957), .CO(n528), .S(n529) );
  CFA1X1 U451 ( .A(n857), .B(n1011), .CI(n911), .CO(n530), .S(n531) );
  CFA1X1 U452 ( .A(n843), .B(n983), .CI(n873), .CO(n532), .S(n533) );
  CFA1X1 U453 ( .A(n813), .B(n831), .CI(n821), .CO(n534), .S(n535) );
  CFA1X1 U454 ( .A(n541), .B(n539), .CI(n560), .CO(n536), .S(n537) );
  CFA1X1 U455 ( .A(n1631), .B(n562), .CI(n543), .CO(n538), .S(n539) );
  CFA1X1 U456 ( .A(n1624), .B(n1626), .CI(n1629), .CO(n540), .S(n541) );
  CFA1X1 U457 ( .A(n1627), .B(n1622), .CI(n1628), .CO(n542), .S(n543) );
  CFA1X1 U458 ( .A(n572), .B(n553), .CI(n555), .CO(n544), .S(n545) );
  CFA1X1 U459 ( .A(n576), .B(n570), .CI(n574), .CO(n546), .S(n547) );
  CFA1X1 U460 ( .A(n912), .B(n557), .CI(n934), .CO(n548), .S(n549) );
  CFA1X1 U461 ( .A(n892), .B(n1042), .CI(n958), .CO(n550), .S(n551) );
  CFA1X1 U462 ( .A(n844), .B(n984), .CI(n858), .CO(n552), .S(n553) );
  CFA1X1 U463 ( .A(n822), .B(n1012), .CI(n874), .CO(n554), .S(n555) );
  CHA1X1 U464 ( .A(n782), .B(n832), .CO(n556), .S(n557) );
  CFA1X1 U465 ( .A(n563), .B(n561), .CI(n580), .CO(n558), .S(n559) );
  CFA1X1 U466 ( .A(n1623), .B(n582), .CI(n1625), .CO(n560), .S(n561) );
  CFA1X1 U467 ( .A(n1618), .B(n1620), .CI(n1621), .CO(n562), .S(n563) );
  CFA1X1 U468 ( .A(n573), .B(n588), .CI(n571), .CO(n564), .S(n565) );
  CFA1X1 U469 ( .A(n590), .B(n575), .CI(n577), .CO(n566), .S(n567) );
  CFA1X1 U470 ( .A(n596), .B(n592), .CI(n594), .CO(n568), .S(n569) );
  CFA1X1 U471 ( .A(n893), .B(n959), .CI(n935), .CO(n570), .S(n571) );
  CFA1X1 U472 ( .A(n875), .B(n1013), .CI(n1043), .CO(n572), .S(n573) );
  CFA1X1 U473 ( .A(n859), .B(n985), .CI(n913), .CO(n574), .S(n575) );
  CFA1X1 U474 ( .A(n823), .B(n845), .CI(n833), .CO(n576), .S(n577) );
  CFA1X1 U475 ( .A(n583), .B(n581), .CI(n600), .CO(n578), .S(n579) );
  CFA1X1 U476 ( .A(n1617), .B(n602), .CI(n1619), .CO(n580), .S(n581) );
  CFA1X1 U477 ( .A(n1613), .B(n1615), .CI(n1616), .CO(n582), .S(n583) );
  CFA1X1 U478 ( .A(n608), .B(n591), .CI(n593), .CO(n584), .S(n585) );
  CFA1X1 U479 ( .A(n610), .B(n595), .CI(n612), .CO(n586), .S(n587) );
  CFA1X1 U480 ( .A(n936), .B(n614), .CI(n597), .CO(n588), .S(n589) );
  CFA1X1 U481 ( .A(n894), .B(n1044), .CI(n960), .CO(n590), .S(n591) );
  CFA1X1 U482 ( .A(n860), .B(n1014), .CI(n914), .CO(n592), .S(n593) );
  CFA1X1 U483 ( .A(n846), .B(n986), .CI(n876), .CO(n594), .S(n595) );
  CHA1X1 U484 ( .A(n783), .B(n834), .CO(n596), .S(n597) );
  CFA1X1 U485 ( .A(n603), .B(n601), .CI(n618), .CO(n598), .S(n599) );
  CFA1X1 U486 ( .A(n1612), .B(n620), .CI(n1614), .CO(n600), .S(n601) );
  CFA1X1 U487 ( .A(n1611), .B(n1610), .CI(n1608), .CO(n602), .S(n603) );
  CFA1X1 U488 ( .A(n615), .B(n611), .CI(n613), .CO(n604), .S(n605) );
  CFA1X1 U489 ( .A(n630), .B(n628), .CI(n626), .CO(n606), .S(n607) );
  CFA1X1 U491 ( .A(n895), .B(n1015), .CI(n961), .CO(n610), .S(n611) );
  CFA1X1 U492 ( .A(n877), .B(n987), .CI(n1045), .CO(n612), .S(n613) );
  CFA1X1 U493 ( .A(n835), .B(n861), .CI(n847), .CO(n614), .S(n615) );
  CFA1X1 U494 ( .A(n621), .B(n619), .CI(n636), .CO(n616), .S(n617) );
  CFA1X1 U495 ( .A(n1607), .B(n638), .CI(n1609), .CO(n618), .S(n619) );
  CFA1X1 U496 ( .A(n1606), .B(n1605), .CI(n1603), .CO(n620), .S(n621) );
  CFA1X1 U497 ( .A(n646), .B(n629), .CI(n631), .CO(n622), .S(n623) );
  CFA1X1 U498 ( .A(n633), .B(n644), .CI(n648), .CO(n624), .S(n625) );
  CFA1X1 U499 ( .A(n916), .B(n962), .CI(n938), .CO(n626), .S(n627) );
  CFA1X1 U500 ( .A(n896), .B(n1016), .CI(n1046), .CO(n628), .S(n629) );
  CFA1X1 U501 ( .A(n848), .B(n988), .CI(n862), .CO(n630), .S(n631) );
  CHA1X1 U502 ( .A(n784), .B(n878), .CO(n632), .S(n633) );
  CFA1X1 U503 ( .A(n639), .B(n637), .CI(n652), .CO(n634), .S(n635) );
  CFA1X1 U504 ( .A(n1602), .B(n1600), .CI(n1604), .CO(n636), .S(n637) );
  CFA1X1 U505 ( .A(n1601), .B(n1598), .CI(n1596), .CO(n638), .S(n639) );
  CFA1X1 U506 ( .A(n660), .B(n647), .CI(n649), .CO(n640), .S(n641) );
  CFA1X1 U507 ( .A(n939), .B(n662), .CI(n664), .CO(n642), .S(n643) );
  CFA1X1 U508 ( .A(n917), .B(n1047), .CI(n963), .CO(n644), .S(n645) );
  CFA1X1 U509 ( .A(n897), .B(n1017), .CI(n989), .CO(n646), .S(n647) );
  CFA1X1 U510 ( .A(n849), .B(n879), .CI(n863), .CO(n648), .S(n649) );
  CFA1X1 U511 ( .A(n1599), .B(n653), .CI(n668), .CO(n650), .S(n651) );
  CFA1X1 U512 ( .A(n1595), .B(n1594), .CI(n1597), .CO(n652), .S(n653) );
  CFA1X1 U513 ( .A(n663), .B(n672), .CI(n661), .CO(n654), .S(n655) );
  CFA1X1 U514 ( .A(n678), .B(n674), .CI(n676), .CO(n656), .S(n657) );
  CFA1X1 U515 ( .A(n898), .B(n665), .CI(n964), .CO(n658), .S(n659) );
  CFA1X1 U516 ( .A(n880), .B(n990), .CI(n1048), .CO(n660), .S(n661) );
  CHA1X1 U518 ( .A(n785), .B(n940), .CO(n664), .S(n665) );
  CFA1X1 U519 ( .A(n1593), .B(n669), .CI(n682), .CO(n666), .S(n667) );
  CFA1X1 U520 ( .A(n1589), .B(n1591), .CI(n1592), .CO(n668), .S(n669) );
  CFA1X1 U521 ( .A(n679), .B(n675), .CI(n677), .CO(n670), .S(n671) );
  CFA1X1 U522 ( .A(n692), .B(n690), .CI(n688), .CO(n672), .S(n673) );
  CFA1X1 U523 ( .A(n941), .B(n1049), .CI(n965), .CO(n674), .S(n675) );
  CFA1X1 U524 ( .A(n919), .B(n1019), .CI(n991), .CO(n676), .S(n677) );
  CFA1X1 U525 ( .A(n865), .B(n899), .CI(n881), .CO(n678), .S(n679) );
  CFA1X1 U526 ( .A(n1590), .B(n683), .CI(n696), .CO(n680), .S(n681) );
  CFA1X1 U527 ( .A(n1585), .B(n1588), .CI(n1587), .CO(n682), .S(n683) );
  CFA1X1 U528 ( .A(n702), .B(n689), .CI(n691), .CO(n684), .S(n685) );
  CFA1X1 U529 ( .A(n920), .B(n704), .CI(n693), .CO(n686), .S(n687) );
  CFA1X1 U530 ( .A(n900), .B(n966), .CI(n942), .CO(n688), .S(n689) );
  CFA1X1 U531 ( .A(n882), .B(n992), .CI(n1050), .CO(n690), .S(n691) );
  CHA1X1 U532 ( .A(n786), .B(n1020), .CO(n692), .S(n693) );
  CFA1X1 U533 ( .A(n1586), .B(n697), .CI(n708), .CO(n694), .S(n695) );
  CFA1X1 U534 ( .A(n1583), .B(n1582), .CI(n1584), .CO(n696), .S(n697) );
  CFA1X1 U535 ( .A(n712), .B(n705), .CI(n714), .CO(n698), .S(n699) );
  CFA1X1 U536 ( .A(n967), .B(n716), .CI(n1051), .CO(n700), .S(n701) );
  CFA1X1 U537 ( .A(n943), .B(n993), .CI(n1021), .CO(n702), .S(n703) );
  CFA1X1 U538 ( .A(n883), .B(n921), .CI(n901), .CO(n704), .S(n705) );
  CFA1X1 U539 ( .A(n1581), .B(n709), .CI(n1578), .CO(n706), .S(n707) );
  CFA1X1 U540 ( .A(n1579), .B(n1576), .CI(n1580), .CO(n708), .S(n709) );
  CFA1X1 U541 ( .A(n717), .B(n724), .CI(n726), .CO(n710), .S(n711) );
  CFA1X1 U542 ( .A(n922), .B(n968), .CI(n944), .CO(n712), .S(n713) );
  CFA1X1 U543 ( .A(n902), .B(n994), .CI(n1052), .CO(n714), .S(n715) );
  CHA1X1 U544 ( .A(n787), .B(n1022), .CO(n716), .S(n717) );
  CFA1X1 U545 ( .A(n1574), .B(n1577), .CI(n1575), .CO(n718), .S(n719) );
  CFA1X1 U546 ( .A(n727), .B(n732), .CI(n725), .CO(n720), .S(n721) );
  CFA1X1 U547 ( .A(n1053), .B(n734), .CI(n736), .CO(n722), .S(n723) );
  CFA1X1 U548 ( .A(n969), .B(n1023), .CI(n995), .CO(n724), .S(n725) );
  CFA1X1 U549 ( .A(n903), .B(n945), .CI(n923), .CO(n726), .S(n727) );
  CFA1X1 U550 ( .A(n1572), .B(n1573), .CI(n1571), .CO(n728), .S(n729) );
  CFA1X1 U551 ( .A(n744), .B(n735), .CI(n742), .CO(n730), .S(n731) );
  CFA1X1 U552 ( .A(n946), .B(n737), .CI(n970), .CO(n732), .S(n733) );
  CFA1X1 U553 ( .A(n924), .B(n996), .CI(n1054), .CO(n734), .S(n735) );
  CHA1X1 U554 ( .A(n788), .B(n1024), .CO(n736), .S(n737) );
  CFA1X1 U555 ( .A(n1569), .B(n1570), .CI(n1566), .CO(n738), .S(n739) );
  CFA1X1 U556 ( .A(n752), .B(n745), .CI(n750), .CO(n740), .S(n741) );
  CFA1X1 U557 ( .A(n1055), .B(n1025), .CI(n997), .CO(n742), .S(n743) );
  CFA1X1 U558 ( .A(n925), .B(n971), .CI(n947), .CO(n744), .S(n745) );
  CFA1X1 U559 ( .A(n756), .B(n749), .CI(n751), .CO(n746), .S(n747) );
  CFA1X1 U560 ( .A(n972), .B(n758), .CI(n753), .CO(n748), .S(n749) );
  CFA1X1 U561 ( .A(n948), .B(n998), .CI(n1056), .CO(n750), .S(n751) );
  CHA1X1 U562 ( .A(n789), .B(n1026), .CO(n752), .S(n753) );
  CFA1X1 U563 ( .A(n762), .B(n757), .CI(n759), .CO(n754), .S(n755) );
  CFA1X1 U564 ( .A(n1027), .B(n764), .CI(n999), .CO(n756), .S(n757) );
  CFA1X1 U565 ( .A(n949), .B(n1057), .CI(n973), .CO(n758), .S(n759) );
  CFA1X1 U566 ( .A(n765), .B(n763), .CI(n768), .CO(n760), .S(n761) );
  CFA1X1 U567 ( .A(n974), .B(n1000), .CI(n1058), .CO(n762), .S(n763) );
  CHA1X1 U568 ( .A(n790), .B(n1028), .CO(n764), .S(n765) );
  CFA1X1 U569 ( .A(n1001), .B(n769), .CI(n772), .CO(n766), .S(n767) );
  CFA1X1 U570 ( .A(n975), .B(n1029), .CI(n1059), .CO(n768), .S(n769) );
  CFA1X1 U571 ( .A(n1030), .B(n773), .CI(n1002), .CO(n770), .S(n771) );
  CHA1X1 U572 ( .A(n1060), .B(n791), .CO(n772), .S(n773) );
  CFA1X1 U573 ( .A(n1003), .B(n1031), .CI(n1061), .CO(n774), .S(n775) );
  CHA1X1 U574 ( .A(n1062), .B(n1032), .CO(n776), .S(n777) );
  COND2X1 U575 ( .A(n115), .B(n1410), .C(n114), .D(n1067), .Z(n778) );
  COND2X1 U576 ( .A(n1065), .B(n114), .C(n115), .D(n1066), .Z(n794) );
  COND2X1 U581 ( .A(n112), .B(n1411), .C(n110), .D(n1072), .Z(n779) );
  COND2X1 U582 ( .A(n1068), .B(n110), .C(n1069), .D(n112), .Z(n796) );
  COND2X1 U583 ( .A(n1070), .B(n112), .C(n110), .D(n1069), .Z(n797) );
  COND2X1 U584 ( .A(n1070), .B(n110), .C(n112), .D(n1071), .Z(n798) );
  COND2X1 U591 ( .A(n107), .B(n1412), .C(n105), .D(n1079), .Z(n780) );
  COND2X1 U592 ( .A(n1073), .B(n105), .C(n1074), .D(n107), .Z(n800) );
  COND2X1 U593 ( .A(n1075), .B(n107), .C(n105), .D(n1074), .Z(n801) );
  COND2X1 U594 ( .A(n1075), .B(n105), .C(n1076), .D(n107), .Z(n802) );
  COND2X1 U595 ( .A(n1077), .B(n107), .C(n105), .D(n1076), .Z(n803) );
  COND2X1 U596 ( .A(n1077), .B(n105), .C(n107), .D(n1078), .Z(n804) );
  CND2IX1 U604 ( .B(n1704), .A(n104), .Z(n1079) );
  COND2X1 U605 ( .A(n102), .B(n1764), .C(n100), .D(n1088), .Z(n781) );
  COND2X1 U607 ( .A(n1082), .B(n102), .C(n1081), .D(n100), .Z(n807) );
  COND2X1 U608 ( .A(n1082), .B(n100), .C(n1083), .D(n102), .Z(n808) );
  COND2X1 U609 ( .A(n1084), .B(n102), .C(n1083), .D(n100), .Z(n809) );
  COND2X1 U610 ( .A(n1084), .B(n100), .C(n1085), .D(n102), .Z(n810) );
  COND2X1 U611 ( .A(n1086), .B(n102), .C(n1085), .D(n100), .Z(n811) );
  COND2X1 U612 ( .A(n1086), .B(n100), .C(n102), .D(n1087), .Z(n812) );
  CND2IX1 U622 ( .B(n1704), .A(n1763), .Z(n1088) );
  COND2X1 U623 ( .A(n97), .B(n1762), .C(n1099), .D(n95), .Z(n782) );
  COND2X1 U624 ( .A(n97), .B(n1090), .C(n95), .D(n1089), .Z(n814) );
  COND2X1 U626 ( .A(n97), .B(n1092), .C(n95), .D(n1091), .Z(n816) );
  COND2X1 U628 ( .A(n1093), .B(n95), .C(n1094), .D(n97), .Z(n818) );
  COND2X1 U630 ( .A(n1095), .B(n95), .C(n1096), .D(n97), .Z(n820) );
  COND2X1 U632 ( .A(n1097), .B(n95), .C(n1098), .D(n97), .Z(n822) );
  CND2IX1 U644 ( .B(n1704), .A(n1761), .Z(n1099) );
  COND2X1 U645 ( .A(n91), .B(n1759), .C(n1112), .D(n89), .Z(n783) );
  COND2X1 U646 ( .A(n91), .B(n1101), .C(n89), .D(n1100), .Z(n824) );
  COND2X1 U647 ( .A(n91), .B(n1102), .C(n1101), .D(n89), .Z(n825) );
  COND2X1 U648 ( .A(n91), .B(n1103), .C(n89), .D(n1102), .Z(n826) );
  COND2X1 U649 ( .A(n91), .B(n1104), .C(n1103), .D(n89), .Z(n827) );
  COND2X1 U650 ( .A(n91), .B(n1105), .C(n89), .D(n1104), .Z(n828) );
  COND2X1 U651 ( .A(n91), .B(n1106), .C(n1105), .D(n89), .Z(n829) );
  COND2X1 U652 ( .A(n91), .B(n1107), .C(n89), .D(n1106), .Z(n830) );
  COND2X1 U653 ( .A(n91), .B(n1108), .C(n1107), .D(n89), .Z(n831) );
  COND2X1 U654 ( .A(n91), .B(n1109), .C(n89), .D(n1108), .Z(n832) );
  COND2X1 U656 ( .A(n91), .B(n1111), .C(n89), .D(n1110), .Z(n834) );
  CND2IX1 U670 ( .B(n1704), .A(n1756), .Z(n1112) );
  COND2X1 U671 ( .A(n84), .B(n1755), .C(n1127), .D(n82), .Z(n784) );
  COND2X1 U672 ( .A(n84), .B(n1114), .C(n1113), .D(n82), .Z(n836) );
  COND2X1 U673 ( .A(n84), .B(n1115), .C(n1114), .D(n82), .Z(n837) );
  COND2X1 U674 ( .A(n84), .B(n1116), .C(n1115), .D(n82), .Z(n838) );
  COND2X1 U675 ( .A(n84), .B(n1117), .C(n1116), .D(n82), .Z(n839) );
  COND2X1 U676 ( .A(n84), .B(n1118), .C(n82), .D(n1117), .Z(n840) );
  COND2X1 U677 ( .A(n84), .B(n1119), .C(n1118), .D(n82), .Z(n841) );
  COND2X1 U678 ( .A(n84), .B(n1120), .C(n82), .D(n1119), .Z(n842) );
  COND2X1 U679 ( .A(n84), .B(n1121), .C(n1120), .D(n82), .Z(n843) );
  COND2X1 U680 ( .A(n84), .B(n1122), .C(n82), .D(n1121), .Z(n844) );
  COND2X1 U681 ( .A(n84), .B(n1123), .C(n1122), .D(n82), .Z(n845) );
  COND2X1 U682 ( .A(n84), .B(n1124), .C(n82), .D(n1123), .Z(n846) );
  COND2X1 U683 ( .A(n84), .B(n1125), .C(n1124), .D(n82), .Z(n847) );
  COND2X1 U684 ( .A(n84), .B(n1126), .C(n82), .D(n1125), .Z(n848) );
  CND2IX1 U700 ( .B(n1704), .A(n1753), .Z(n1127) );
  CND2IX1 U734 ( .B(n1704), .A(n1747), .Z(n1144) );
  COND2X1 U735 ( .A(n69), .B(n1524), .C(n1163), .D(n66), .Z(n786) );
  COND2X1 U736 ( .A(n69), .B(n1146), .C(n1145), .D(n66), .Z(n866) );
  COND2X1 U737 ( .A(n69), .B(n1147), .C(n1146), .D(n66), .Z(n867) );
  COND2X1 U738 ( .A(n69), .B(n1148), .C(n1147), .D(n66), .Z(n868) );
  COND2X1 U739 ( .A(n69), .B(n1149), .C(n1148), .D(n66), .Z(n869) );
  COND2X1 U740 ( .A(n69), .B(n1150), .C(n1149), .D(n66), .Z(n870) );
  COND2X1 U741 ( .A(n69), .B(n1151), .C(n1150), .D(n66), .Z(n871) );
  COND2X1 U742 ( .A(n69), .B(n1152), .C(n1151), .D(n66), .Z(n872) );
  COND2X1 U743 ( .A(n69), .B(n1153), .C(n1152), .D(n66), .Z(n873) );
  COND2X1 U744 ( .A(n69), .B(n1154), .C(n1153), .D(n66), .Z(n874) );
  COND2X1 U745 ( .A(n69), .B(n1155), .C(n1154), .D(n66), .Z(n875) );
  COND2X1 U746 ( .A(n69), .B(n1156), .C(n1155), .D(n66), .Z(n876) );
  COND2X1 U747 ( .A(n69), .B(n1157), .C(n1156), .D(n66), .Z(n877) );
  COND2X1 U748 ( .A(n69), .B(n1158), .C(n66), .D(n1157), .Z(n878) );
  COND2X1 U749 ( .A(n69), .B(n1159), .C(n1158), .D(n66), .Z(n879) );
  COND2X1 U750 ( .A(n69), .B(n1160), .C(n66), .D(n1159), .Z(n880) );
  COND2X1 U752 ( .A(n69), .B(n1162), .C(n66), .D(n1161), .Z(n882) );
  CND2IX1 U772 ( .B(n1704), .A(n1744), .Z(n1163) );
  COND2X1 U790 ( .A(n61), .B(n1181), .C(n58), .D(n1180), .Z(n900) );
  COND2X1 U816 ( .A(n53), .B(n1186), .C(n1185), .D(n50), .Z(n904) );
  COND2X1 U817 ( .A(n53), .B(n1187), .C(n1186), .D(n50), .Z(n905) );
  COND2X1 U818 ( .A(n53), .B(n1188), .C(n1187), .D(n50), .Z(n906) );
  COND2X1 U819 ( .A(n53), .B(n1189), .C(n1188), .D(n50), .Z(n907) );
  COND2X1 U820 ( .A(n53), .B(n1190), .C(n1189), .D(n50), .Z(n908) );
  COND2X1 U821 ( .A(n53), .B(n1191), .C(n1190), .D(n50), .Z(n909) );
  COND2X1 U822 ( .A(n53), .B(n1192), .C(n1191), .D(n50), .Z(n910) );
  COND2X1 U823 ( .A(n53), .B(n1193), .C(n1192), .D(n50), .Z(n911) );
  COND2X1 U824 ( .A(n53), .B(n1194), .C(n1193), .D(n50), .Z(n912) );
  COND2X1 U825 ( .A(n53), .B(n1195), .C(n1194), .D(n50), .Z(n913) );
  COND2X1 U826 ( .A(n53), .B(n1196), .C(n1195), .D(n50), .Z(n914) );
  COND2X1 U827 ( .A(n53), .B(n1197), .C(n1196), .D(n50), .Z(n915) );
  COND2X1 U828 ( .A(n53), .B(n1198), .C(n1197), .D(n50), .Z(n916) );
  COND2X1 U829 ( .A(n53), .B(n1199), .C(n1198), .D(n50), .Z(n917) );
  COND2X1 U830 ( .A(n53), .B(n1200), .C(n1199), .D(n50), .Z(n918) );
  COND2X1 U831 ( .A(n53), .B(n1201), .C(n1200), .D(n50), .Z(n919) );
  COND2X1 U832 ( .A(n53), .B(n1202), .C(n50), .D(n1201), .Z(n920) );
  COND2X1 U834 ( .A(n53), .B(n1204), .C(n50), .D(n1203), .Z(n922) );
  COND2X1 U835 ( .A(n53), .B(n1205), .C(n1204), .D(n50), .Z(n923) );
  COND2X1 U836 ( .A(n53), .B(n1206), .C(n50), .D(n1205), .Z(n924) );
  CND2IX1 U860 ( .B(n1704), .A(n1741), .Z(n1207) );
  COND2X1 U861 ( .A(n44), .B(n1738), .C(n1232), .D(n42), .Z(n789) );
  COND2X1 U862 ( .A(n44), .B(n1209), .C(n1208), .D(n42), .Z(n926) );
  COND2X1 U863 ( .A(n44), .B(n1210), .C(n1209), .D(n42), .Z(n927) );
  COND2X1 U864 ( .A(n44), .B(n1211), .C(n1210), .D(n42), .Z(n928) );
  COND2X1 U865 ( .A(n44), .B(n1212), .C(n1211), .D(n42), .Z(n929) );
  COND2X1 U866 ( .A(n44), .B(n1213), .C(n1212), .D(n42), .Z(n930) );
  COND2X1 U867 ( .A(n44), .B(n1214), .C(n1213), .D(n42), .Z(n931) );
  COND2X1 U868 ( .A(n44), .B(n1215), .C(n1214), .D(n42), .Z(n932) );
  COND2X1 U869 ( .A(n44), .B(n1216), .C(n1215), .D(n42), .Z(n933) );
  COND2X1 U870 ( .A(n44), .B(n1217), .C(n1216), .D(n42), .Z(n934) );
  COND2X1 U871 ( .A(n44), .B(n1218), .C(n1217), .D(n42), .Z(n935) );
  COND2X1 U872 ( .A(n44), .B(n1219), .C(n1218), .D(n42), .Z(n936) );
  COND2X1 U873 ( .A(n44), .B(n1220), .C(n1219), .D(n42), .Z(n937) );
  COND2X1 U874 ( .A(n44), .B(n1221), .C(n1220), .D(n42), .Z(n938) );
  COND2X1 U875 ( .A(n44), .B(n1222), .C(n1221), .D(n42), .Z(n939) );
  COND2X1 U876 ( .A(n44), .B(n1223), .C(n1222), .D(n42), .Z(n940) );
  COND2X1 U877 ( .A(n44), .B(n1224), .C(n1223), .D(n42), .Z(n941) );
  COND2X1 U878 ( .A(n44), .B(n1225), .C(n1224), .D(n42), .Z(n942) );
  COND2X1 U879 ( .A(n44), .B(n1226), .C(n1225), .D(n42), .Z(n943) );
  COND2X1 U880 ( .A(n44), .B(n1227), .C(n1226), .D(n42), .Z(n944) );
  COND2X1 U881 ( .A(n44), .B(n1228), .C(n1227), .D(n42), .Z(n945) );
  COND2X1 U882 ( .A(n44), .B(n1229), .C(n42), .D(n1228), .Z(n946) );
  COND2X1 U883 ( .A(n44), .B(n1230), .C(n1229), .D(n42), .Z(n947) );
  COND2X1 U884 ( .A(n44), .B(n1231), .C(n42), .D(n1230), .Z(n948) );
  CND2IX1 U910 ( .B(n1704), .A(n1736), .Z(n1232) );
  CND2IX1 U964 ( .B(n1704), .A(n1724), .Z(n1259) );
  COND2X1 U965 ( .A(n27), .B(n1723), .C(n1288), .D(n24), .Z(n791) );
  COND2X1 U966 ( .A(n27), .B(n1261), .C(n24), .D(n1260), .Z(n976) );
  COND2X1 U967 ( .A(n27), .B(n1262), .C(n24), .D(n1261), .Z(n977) );
  COND2X1 U968 ( .A(n27), .B(n1263), .C(n24), .D(n1262), .Z(n978) );
  COND2X1 U969 ( .A(n27), .B(n1264), .C(n24), .D(n1263), .Z(n979) );
  COND2X1 U970 ( .A(n27), .B(n1265), .C(n24), .D(n1264), .Z(n980) );
  COND2X1 U971 ( .A(n27), .B(n1266), .C(n24), .D(n1265), .Z(n981) );
  COND2X1 U972 ( .A(n27), .B(n1267), .C(n24), .D(n1266), .Z(n982) );
  COND2X1 U973 ( .A(n27), .B(n1268), .C(n24), .D(n1267), .Z(n983) );
  COND2X1 U974 ( .A(n27), .B(n1269), .C(n24), .D(n1268), .Z(n984) );
  COND2X1 U975 ( .A(n27), .B(n1270), .C(n24), .D(n1269), .Z(n985) );
  COND2X1 U976 ( .A(n27), .B(n1271), .C(n24), .D(n1270), .Z(n986) );
  COND2X1 U977 ( .A(n27), .B(n1272), .C(n24), .D(n1271), .Z(n987) );
  COND2X1 U978 ( .A(n27), .B(n1273), .C(n24), .D(n1272), .Z(n988) );
  COND2X1 U979 ( .A(n27), .B(n1274), .C(n24), .D(n1273), .Z(n989) );
  COND2X1 U980 ( .A(n27), .B(n1275), .C(n24), .D(n1274), .Z(n990) );
  COND2X1 U981 ( .A(n27), .B(n1276), .C(n24), .D(n1275), .Z(n991) );
  COND2X1 U982 ( .A(n27), .B(n1277), .C(n24), .D(n1276), .Z(n992) );
  COND2X1 U983 ( .A(n27), .B(n1278), .C(n24), .D(n1277), .Z(n993) );
  COND2X1 U984 ( .A(n27), .B(n1279), .C(n24), .D(n1278), .Z(n994) );
  COND2X1 U985 ( .A(n27), .B(n1280), .C(n24), .D(n1279), .Z(n995) );
  COND2X1 U986 ( .A(n27), .B(n1281), .C(n24), .D(n1280), .Z(n996) );
  COND2X1 U987 ( .A(n27), .B(n1282), .C(n24), .D(n1281), .Z(n997) );
  COND2X1 U988 ( .A(n27), .B(n1283), .C(n24), .D(n1282), .Z(n998) );
  COND2X1 U989 ( .A(n27), .B(n1284), .C(n24), .D(n1283), .Z(n999) );
  COND2X1 U990 ( .A(n27), .B(n1285), .C(n24), .D(n1284), .Z(n1000) );
  COND2X1 U991 ( .A(n27), .B(n1286), .C(n24), .D(n1285), .Z(n1001) );
  COND2X1 U992 ( .A(n27), .B(n1287), .C(n24), .D(n1286), .Z(n1002) );
  CND2IX1 U1022 ( .B(n1704), .A(n1721), .Z(n1288) );
  COND2X1 U1023 ( .A(n18), .B(n1717), .C(n1319), .D(n15), .Z(n792) );
  COND2X1 U1024 ( .A(n18), .B(n1290), .C(n15), .D(n1289), .Z(n1004) );
  COND2X1 U1025 ( .A(n18), .B(n1291), .C(n15), .D(n1290), .Z(n1005) );
  COND2X1 U1026 ( .A(n18), .B(n1292), .C(n15), .D(n1291), .Z(n1006) );
  COND2X1 U1027 ( .A(n18), .B(n1293), .C(n15), .D(n1292), .Z(n1007) );
  COND2X1 U1028 ( .A(n18), .B(n1294), .C(n15), .D(n1293), .Z(n1008) );
  COND2X1 U1029 ( .A(n18), .B(n1295), .C(n15), .D(n1294), .Z(n1009) );
  COND2X1 U1030 ( .A(n18), .B(n1296), .C(n15), .D(n1295), .Z(n1010) );
  COND2X1 U1031 ( .A(n18), .B(n1297), .C(n15), .D(n1296), .Z(n1011) );
  COND2X1 U1032 ( .A(n18), .B(n1298), .C(n15), .D(n1297), .Z(n1012) );
  COND2X1 U1033 ( .A(n18), .B(n1299), .C(n15), .D(n1298), .Z(n1013) );
  COND2X1 U1034 ( .A(n18), .B(n1300), .C(n15), .D(n1299), .Z(n1014) );
  COND2X1 U1035 ( .A(n18), .B(n1301), .C(n15), .D(n1300), .Z(n1015) );
  COND2X1 U1036 ( .A(n18), .B(n1302), .C(n15), .D(n1301), .Z(n1016) );
  COND2X1 U1037 ( .A(n18), .B(n1303), .C(n15), .D(n1302), .Z(n1017) );
  COND2X1 U1038 ( .A(n18), .B(n1304), .C(n15), .D(n1303), .Z(n1018) );
  COND2X1 U1039 ( .A(n18), .B(n1305), .C(n15), .D(n1304), .Z(n1019) );
  COND2X1 U1040 ( .A(n18), .B(n1306), .C(n15), .D(n1305), .Z(n1020) );
  COND2X1 U1041 ( .A(n18), .B(n1307), .C(n15), .D(n1306), .Z(n1021) );
  COND2X1 U1042 ( .A(n18), .B(n1308), .C(n15), .D(n1307), .Z(n1022) );
  COND2X1 U1043 ( .A(n18), .B(n1309), .C(n15), .D(n1308), .Z(n1023) );
  COND2X1 U1044 ( .A(n18), .B(n1310), .C(n15), .D(n1309), .Z(n1024) );
  COND2X1 U1045 ( .A(n18), .B(n1311), .C(n15), .D(n1310), .Z(n1025) );
  COND2X1 U1046 ( .A(n18), .B(n1312), .C(n15), .D(n1311), .Z(n1026) );
  COND2X1 U1047 ( .A(n18), .B(n1313), .C(n15), .D(n1312), .Z(n1027) );
  COND2X1 U1048 ( .A(n18), .B(n1314), .C(n15), .D(n1313), .Z(n1028) );
  COND2X1 U1050 ( .A(n18), .B(n1316), .C(n15), .D(n1315), .Z(n1030) );
  COND2X1 U1051 ( .A(n18), .B(n1317), .C(n15), .D(n1316), .Z(n1031) );
  COND2X1 U1052 ( .A(n18), .B(n1318), .C(n15), .D(n1317), .Z(n1032) );
  CND2IX1 U1084 ( .B(n1704), .A(n1711), .Z(n1319) );
  COND2X1 U1085 ( .A(n9), .B(n1528), .C(n6), .D(n1352), .Z(n793) );
  COND2X1 U1086 ( .A(n9), .B(n1321), .C(n6), .D(n1320), .Z(n1034) );
  COND2X1 U1087 ( .A(n9), .B(n1322), .C(n6), .D(n1321), .Z(n1035) );
  COND2X1 U1088 ( .A(n9), .B(n1323), .C(n6), .D(n1322), .Z(n1036) );
  COND2X1 U1089 ( .A(n9), .B(n1324), .C(n6), .D(n1323), .Z(n1037) );
  COND2X1 U1090 ( .A(n9), .B(n1325), .C(n6), .D(n1324), .Z(n1038) );
  COND2X1 U1091 ( .A(n9), .B(n1326), .C(n6), .D(n1325), .Z(n1039) );
  COND2X1 U1092 ( .A(n9), .B(n1327), .C(n6), .D(n1326), .Z(n1040) );
  COND2X1 U1093 ( .A(n9), .B(n1328), .C(n6), .D(n1327), .Z(n1041) );
  COND2X1 U1094 ( .A(n9), .B(n1329), .C(n6), .D(n1328), .Z(n1042) );
  COND2X1 U1095 ( .A(n9), .B(n1330), .C(n6), .D(n1329), .Z(n1043) );
  COND2X1 U1096 ( .A(n9), .B(n1331), .C(n6), .D(n1330), .Z(n1044) );
  COND2X1 U1097 ( .A(n9), .B(n1332), .C(n6), .D(n1331), .Z(n1045) );
  COND2X1 U1098 ( .A(n9), .B(n1333), .C(n6), .D(n1332), .Z(n1046) );
  COND2X1 U1099 ( .A(n9), .B(n1334), .C(n6), .D(n1333), .Z(n1047) );
  COND2X1 U1100 ( .A(n9), .B(n1335), .C(n6), .D(n1334), .Z(n1048) );
  COND2X1 U1101 ( .A(n9), .B(n1336), .C(n6), .D(n1335), .Z(n1049) );
  COND2X1 U1102 ( .A(n9), .B(n1337), .C(n6), .D(n1336), .Z(n1050) );
  COND2X1 U1103 ( .A(n9), .B(n1338), .C(n6), .D(n1337), .Z(n1051) );
  COND2X1 U1104 ( .A(n9), .B(n1339), .C(n6), .D(n1338), .Z(n1052) );
  COND2X1 U1105 ( .A(n9), .B(n1340), .C(n6), .D(n1339), .Z(n1053) );
  COND2X1 U1106 ( .A(n9), .B(n1341), .C(n6), .D(n1340), .Z(n1054) );
  COND2X1 U1107 ( .A(n9), .B(n1342), .C(n6), .D(n1341), .Z(n1055) );
  COND2X1 U1108 ( .A(n9), .B(n1343), .C(n6), .D(n1342), .Z(n1056) );
  COND2X1 U1109 ( .A(n9), .B(n1344), .C(n6), .D(n1343), .Z(n1057) );
  COND2X1 U1110 ( .A(n9), .B(n1345), .C(n6), .D(n1344), .Z(n1058) );
  COND2X1 U1111 ( .A(n9), .B(n1346), .C(n6), .D(n1345), .Z(n1059) );
  COND2X1 U1113 ( .A(n9), .B(n1348), .C(n6), .D(n1347), .Z(n1061) );
  COND2X1 U1114 ( .A(n9), .B(n1349), .C(n6), .D(n1348), .Z(n1062) );
  COND2X1 U1115 ( .A(n9), .B(n1350), .C(n6), .D(n1349), .Z(n1063) );
  COND2X1 U1116 ( .A(n9), .B(n1351), .C(n6), .D(n1350), .Z(n1064) );
  CENX2 U1228 ( .A(n1734), .B(a[10]), .Z(n50) );
  CFD1QXL clk_r_REG8_S1 ( .D(n348), .CP(n1692), .Q(n1684) );
  CFD1QXL clk_r_REG2_S1 ( .D(n370), .CP(n1692), .Q(n1678) );
  CFD1QXL clk_r_REG4_S1 ( .D(n350), .CP(n1692), .Q(n1682) );
  CFD1QXL clk_r_REG3_S1 ( .D(n371), .CP(n1692), .Q(n1677) );
  CFD1QXL clk_r_REG7_S1 ( .D(n375), .CP(n1692), .Q(n1674) );
  CFD1QXL clk_r_REG17_S1 ( .D(n399), .CP(n1692), .Q(n1670) );
  CFD1QXL clk_r_REG32_S1 ( .D(n475), .CP(n1692), .Q(n1650) );
  CFD1QXL clk_r_REG58_S1 ( .D(n453), .CP(n1692), .Q(n1656) );
  CFD1QXL clk_r_REG13_S1 ( .D(n427), .CP(n1692), .Q(n1663) );
  CFD1QXL clk_r_REG60_S1 ( .D(n499), .CP(n1692), .Q(n1644) );
  CFD1QXL clk_r_REG39_S1 ( .D(n523), .CP(n1692), .Q(n1638) );
  CFD1QXL clk_r_REG30_S1 ( .D(n503), .CP(n1692), .Q(n1640) );
  CFD1QXL clk_r_REG45_S1 ( .D(n479), .CP(n1692), .Q(n1646) );
  CFD1QXL clk_r_REG80_S1 ( .D(n654), .CP(n1692), .Q(n1600) );
  CFD1QXL clk_r_REG101_S1 ( .D(n721), .CP(n1692), .Q(n1577) );
  CFD1QXL clk_r_REG107_S1 ( .D(n731), .CP(n1692), .Q(n1573) );
  CFD1QXL clk_r_REG70_S1 ( .D(n622), .CP(n1692), .Q(n1610) );
  CFD1QXL clk_r_REG66_S1 ( .D(n584), .CP(n1692), .Q(n1620) );
  CFD1QXL clk_r_REG82_S1 ( .D(n670), .CP(n1692), .Q(n1594) );
  CFD1QXL clk_r_REG84_S1 ( .D(n656), .CP(n1692), .Q(n1598) );
  CFD1QXL clk_r_REG112_S1 ( .D(n741), .CP(n1692), .Q(n1570) );
  CFD1QXL clk_r_REG89_S1 ( .D(n684), .CP(n1692), .Q(n1591) );
  CFD1QXL clk_r_REG87_S1 ( .D(n687), .CP(n1692), .Q(n1588) );
  CFD1QXL clk_r_REG103_S1 ( .D(n722), .CP(n1692), .Q(n1576) );
  CFD1QXL clk_r_REG1_S1 ( .D(n351), .CP(n1692), .Q(n1681) );
  CFD1QXL clk_r_REG10_S1 ( .D(n368), .CP(n1692), .Q(n1680) );
  CFD1QXL clk_r_REG122_S1 ( .D(n287), .CP(n1692), .Q(n1688) );
  CFD1QXL clk_r_REG124_S1 ( .D(n1557), .CP(n1692), .Q(n1690) );
  CFD1QXL clk_r_REG120_S1 ( .D(n1545), .CP(n1692), .Q(n1691) );
  CFD1QXL clk_r_REG121_S1 ( .D(n288), .CP(n1692), .Q(n1687) );
  CFD1QXL clk_r_REG28_S1 ( .D(n477), .CP(n1692), .Q(n1648) );
  CFD1QXL clk_r_REG116_S1 ( .D(n457), .CP(n1692), .Q(n1653) );
  CFD1QXL clk_r_REG27_S1 ( .D(n476), .CP(n1692), .Q(n1649) );
  CFD1QXL clk_r_REG20_S1 ( .D(n424), .CP(n1692), .Q(n1666) );
  CFD1QXL clk_r_REG23_S1 ( .D(n428), .CP(n1692), .Q(n1662) );
  CFD1QXL clk_r_REG33_S1 ( .D(n450), .CP(n1692), .Q(n1659) );
  CFD1QXL clk_r_REG34_S1 ( .D(n451), .CP(n1692), .Q(n1658) );
  CFD1QXL clk_r_REG25_S1 ( .D(n454), .CP(n1692), .Q(n1655) );
  CFD1QXL clk_r_REG43_S1 ( .D(n501), .CP(n1692), .Q(n1642) );
  CFD1QXL clk_r_REG36_S1 ( .D(n525), .CP(n1692), .Q(n1636) );
  CFD1QXL clk_r_REG35_S1 ( .D(n524), .CP(n1692), .Q(n1637) );
  CFD1QXL clk_r_REG42_S1 ( .D(n500), .CP(n1692), .Q(n1643) );
  CFD1QXL clk_r_REG75_S1 ( .D(n641), .CP(n1692), .Q(n1604) );
  CFD1QXL clk_r_REG62_S1 ( .D(n605), .CP(n1692), .Q(n1614) );
  CFD1QXL clk_r_REG67_S1 ( .D(n585), .CP(n1692), .Q(n1619) );
  CFD1QXL clk_r_REG71_S1 ( .D(n623), .CP(n1692), .Q(n1609) );
  CFD1QXL clk_r_REG54_S1 ( .D(n565), .CP(n1692), .Q(n1625) );
  CFD1QXL clk_r_REG100_S1 ( .D(n720), .CP(n1692), .Q(n1578) );
  CFD1QXL clk_r_REG113_S1 ( .D(n748), .CP(n1692), .Q(n1566) );
  CFD1QXL clk_r_REG88_S1 ( .D(n673), .CP(n1692), .Q(n1592) );
  CFD1QXL clk_r_REG11_S1 ( .D(n369), .CP(n1692), .Q(n1679) );
  CFD1QXL clk_r_REG5_S1 ( .D(n396), .CP(n1692), .Q(n1673) );
  CFD1QXL clk_r_REG6_S1 ( .D(n397), .CP(n1692), .Q(n1672) );
  CFD1QXL clk_r_REG14_S1 ( .D(n400), .CP(n1692), .Q(n1669) );
  CFD1QXL clk_r_REG21_S1 ( .D(n425), .CP(n1692), .Q(n1665) );
  CFD1QXL clk_r_REG59_S1 ( .D(n498), .CP(n1692), .Q(n1645) );
  CFD1QXL clk_r_REG22_S1 ( .D(n463), .CP(n1692), .Q(n1652) );
  CFD1QXL clk_r_REG26_S1 ( .D(n455), .CP(n1692), .Q(n1654) );
  CFD1QXL clk_r_REG9_S1 ( .D(n403), .CP(n1692), .Q(n1667) );
  CFD1QXL clk_r_REG105_S1 ( .D(n431), .CP(n1692), .Q(n1660) );
  CFD1QXL clk_r_REG31_S1 ( .D(n474), .CP(n1692), .Q(n1651) );
  CFD1QXL clk_r_REG38_S1 ( .D(n522), .CP(n1692), .Q(n1639) );
  CFD1QXL clk_r_REG46_S1 ( .D(n544), .CP(n1692), .Q(n1632) );
  CFD1QXL clk_r_REG29_S1 ( .D(n502), .CP(n1692), .Q(n1641) );
  CFD1QXL clk_r_REG40_S1 ( .D(n526), .CP(n1692), .Q(n1635) );
  CFD1QXL clk_r_REG81_S1 ( .D(n655), .CP(n1692), .Q(n1599) );
  CFD1QXL clk_r_REG79_S1 ( .D(n643), .CP(n1692), .Q(n1602) );
  CFD1QXL clk_r_REG106_S1 ( .D(n730), .CP(n1692), .Q(n1574) );
  CFD1QXL clk_r_REG92_S1 ( .D(n699), .CP(n1692), .Q(n1586) );
  CFD1QXL clk_r_REG83_S1 ( .D(n671), .CP(n1692), .Q(n1593) );
  CFD1QXL clk_r_REG47_S1 ( .D(n545), .CP(n1692), .Q(n1631) );
  CFD1QXL clk_r_REG73_S1 ( .D(n607), .CP(n1692), .Q(n1612) );
  CFD1QXL clk_r_REG69_S1 ( .D(n587), .CP(n1692), .Q(n1617) );
  CFD1QXL clk_r_REG49_S1 ( .D(n567), .CP(n1692), .Q(n1623) );
  CFD1QXL clk_r_REG127_S1 ( .D(n743), .CP(n1692), .Q(n1569) );
  CFD1QXL clk_r_REG94_S1 ( .D(n711), .CP(n1692), .Q(n1581) );
  CFD1QXL clk_r_REG119_S1 ( .D(n285), .CP(n1692), .Q(n1689) );
  CFD1QXL clk_r_REG123_S1 ( .D(n293), .CP(n1692), .Q(n1686) );
  CFD1QXL clk_r_REG115_S1 ( .D(n747), .CP(n1692), .Q(n1567) );
  CFD1QXL clk_r_REG126_S1 ( .D(n294), .CP(n1692), .Q(n1685) );
  CFD1QX1 clk_r_REG98_S1 ( .D(n715), .CP(n1692), .Q(n1579) );
  CFD1QX1 clk_r_REG99_S1 ( .D(n551), .CP(n1692), .Q(n1627) );
  CFD1QX2 clk_r_REG117_S1 ( .D(n703), .CP(n1692), .Q(n1583) );
  CFD1QX1 clk_r_REG97_S1 ( .D(n529), .CP(n1692), .Q(n1633) );
  CFD1QX1 clk_r_REG72_S1 ( .D(n606), .CP(n1692), .Q(n1613) );
  CFD1QX1 clk_r_REG110_S1 ( .D(n627), .CP(n1692), .Q(n1606) );
  CFD1QX1 clk_r_REG78_S1 ( .D(n642), .CP(n1692), .Q(n1603) );
  CFD1QX1 clk_r_REG50_S1 ( .D(n546), .CP(n1692), .Q(n1630) );
  CFD1QX2 clk_r_REG77_S1 ( .D(n659), .CP(n1692), .Q(n1595) );
  CFD1QX1 clk_r_REG37_S1 ( .D(n549), .CP(n1692), .Q(n1628) );
  CFD1QX1 clk_r_REG55_S1 ( .D(n568), .CP(n1692), .Q(n1622) );
  CFD1QX1 clk_r_REG96_S1 ( .D(n701), .CP(n1692), .Q(n1584) );
  CFD1QX1 clk_r_REG48_S1 ( .D(n566), .CP(n1692), .Q(n1624) );
  CFD1QX1 clk_r_REG86_S1 ( .D(n686), .CP(n1692), .Q(n1589) );
  CFD1QX2 clk_r_REG51_S1 ( .D(n547), .CP(n1692), .Q(n1629) );
  CFD1QX1 clk_r_REG41_S1 ( .D(n527), .CP(n1692), .Q(n1634) );
  CFD1QX1 clk_r_REG52_S1 ( .D(n589), .CP(n1692), .Q(n1616) );
  CFD1QXL clk_r_REG18_S1 ( .D(n372), .CP(n1692), .Q(n1676) );
  CFD1QXL clk_r_REG0_S1 ( .D(n349), .CP(n1692), .Q(n1683) );
  CFD1QXL clk_r_REG102_S1 ( .D(n733), .CP(n1692), .Q(n1572) );
  CFD1QXL clk_r_REG44_S1 ( .D(n478), .CP(n1692), .Q(n1647) );
  CFD1QXL clk_r_REG118_S1 ( .D(n754), .CP(n1692), .Q(n1565) );
  CFD1QXL clk_r_REG111_S1 ( .D(n740), .CP(n1692), .Q(n1571) );
  CFD1QXL clk_r_REG57_S1 ( .D(n452), .CP(n1692), .Q(n1657) );
  CFD1QXL clk_r_REG15_S1 ( .D(n401), .CP(n1692), .Q(n1668) );
  CFD1QXL clk_r_REG12_S1 ( .D(n426), .CP(n1692), .Q(n1664) );
  CFD1QXL clk_r_REG24_S1 ( .D(n429), .CP(n1692), .Q(n1661) );
  CFD1QXL clk_r_REG16_S1 ( .D(n398), .CP(n1692), .Q(n1671) );
  CFD1QXL clk_r_REG90_S1 ( .D(n685), .CP(n1692), .Q(n1590) );
  CFD1QXL clk_r_REG104_S1 ( .D(n723), .CP(n1692), .Q(n1575) );
  CFD1QXL clk_r_REG19_S1 ( .D(n373), .CP(n1692), .Q(n1675) );
  CFD1QXL clk_r_REG64_S1 ( .D(n625), .CP(n1692), .Q(n1607) );
  CFD1QXL clk_r_REG114_S1 ( .D(n746), .CP(n1692), .Q(n1568) );
  CFD1QX1 clk_r_REG85_S1 ( .D(n657), .CP(n1692), .Q(n1597) );
  CFD1QX2 clk_r_REG65_S1 ( .D(n609), .CP(n1692), .Q(n1611) );
  CFD1QX1 clk_r_REG53_S1 ( .D(n564), .CP(n1692), .Q(n1626) );
  CFD1QX1 clk_r_REG109_S1 ( .D(n645), .CP(n1692), .Q(n1601) );
  CFD1QX1 clk_r_REG68_S1 ( .D(n586), .CP(n1692), .Q(n1618) );
  CFD1QX1 clk_r_REG63_S1 ( .D(n624), .CP(n1692), .Q(n1608) );
  CFD1QX1 clk_r_REG76_S1 ( .D(n658), .CP(n1692), .Q(n1596) );
  CFD1QX1 clk_r_REG56_S1 ( .D(n569), .CP(n1692), .Q(n1621) );
  CFD1QX1 clk_r_REG61_S1 ( .D(n604), .CP(n1692), .Q(n1615) );
  CFD1QX1 clk_r_REG95_S1 ( .D(n700), .CP(n1692), .Q(n1585) );
  CFD1QX1 clk_r_REG93_S1 ( .D(n710), .CP(n1692), .Q(n1582) );
  CFD1QX1 clk_r_REG108_S1 ( .D(n713), .CP(n1692), .Q(n1580) );
  CFD1QX1 clk_r_REG91_S1 ( .D(n698), .CP(n1692), .Q(n1587) );
  CFD1QX1 clk_r_REG74_S1 ( .D(n640), .CP(n1692), .Q(n1605) );
  CANR1X2 U1246 ( .A(n217), .B(n1550), .C(n212), .Z(n210) );
  CANR1X1 U1247 ( .A(n241), .B(n222), .C(n223), .Z(n221) );
  CIVX2 U1248 ( .A(n1563), .Z(n33) );
  CDLY1XL U1249 ( .A(n1383), .Z(n1706) );
  CNIVX1 U1250 ( .A(n1380), .Z(n1694) );
  CENX1 U1251 ( .A(n1721), .B(n1694), .Z(n1283) );
  CENX1 U1252 ( .A(n1705), .B(n1741), .Z(n1205) );
  CENX1 U1253 ( .A(n1715), .B(n1700), .Z(n1308) );
  CENX1 U1254 ( .A(n1753), .B(n1696), .Z(n1120) );
  CENX1 U1255 ( .A(n1694), .B(n104), .Z(n1074) );
  CANR1X1 U1256 ( .A(n1558), .B(n250), .C(n245), .Z(n243) );
  CENX1 U1257 ( .A(n1740), .B(n1700), .Z(n1196) );
  CENX1 U1258 ( .A(n1721), .B(n1700), .Z(n1277) );
  CENX1 U1259 ( .A(n1735), .B(n1700), .Z(n1221) );
  COND2XL U1260 ( .A(n36), .B(n1250), .C(n1249), .D(n33), .Z(n966) );
  CIVDXL U1261 ( .A(n79), .Z0(n1522), .Z1(n1523) );
  CIVX1 U1262 ( .A(n1524), .Z(n1745) );
  CIVX1 U1263 ( .A(n1524), .Z(n1746) );
  CIVX2 U1264 ( .A(n1524), .Z(n1744) );
  CIVX1 U1265 ( .A(n39), .Z(n1739) );
  CIVDXL U1266 ( .A(n63), .Z0(n1524), .Z1(n1525) );
  CIVX1 U1267 ( .A(n1717), .Z(n1712) );
  CIVDXL U1268 ( .A(n55), .Z0(n1526), .Z1(n1527) );
  CIVDX1 U1269 ( .A(n3), .Z0(n1528), .Z1(n1529) );
  CAN2X1 U1270 ( .A(n1541), .B(n312), .Z(product[1]) );
  CFA1XL U1271 ( .A(n830), .B(n890), .CI(n856), .CO(n508), .S(n509) );
  CFA1XL U1272 ( .A(n855), .B(n1009), .CI(n909), .CO(n484), .S(n485) );
  CFA1XL U1273 ( .A(n864), .B(n1018), .CI(n918), .CO(n662), .S(n663) );
  COND1X1 U1274 ( .A(n257), .B(n251), .C(n252), .Z(n250) );
  COND1X1 U1275 ( .A(n167), .B(n1535), .C(n168), .Z(n166) );
  CANR1X1 U1276 ( .A(n175), .B(n1552), .C(n170), .Z(n168) );
  CEOX1 U1277 ( .A(a[2]), .B(n1712), .Z(n1399) );
  CFA1X2 U1278 ( .A(n915), .B(n632), .CI(n937), .CO(n608), .S(n609) );
  CENX2 U1279 ( .A(n1748), .B(a[18]), .Z(n82) );
  CND2X4 U1280 ( .A(n1391), .B(n82), .Z(n84) );
  CANR1X1 U1281 ( .A(n237), .B(n1559), .C(n230), .Z(n228) );
  CIVX1 U1282 ( .A(n235), .Z(n237) );
  CEOX1 U1283 ( .A(a[10]), .B(n1741), .Z(n1395) );
  CIVX2 U1284 ( .A(n1742), .Z(n1741) );
  CENXL U1285 ( .A(n1741), .B(n1368), .Z(n1190) );
  CENXL U1286 ( .A(n1741), .B(n1370), .Z(n1192) );
  CENXL U1287 ( .A(n1741), .B(n1372), .Z(n1194) );
  CENXL U1288 ( .A(n1695), .B(n1741), .Z(n1201) );
  COND2XL U1289 ( .A(n53), .B(n1742), .C(n1207), .D(n50), .Z(n788) );
  CND2IX4 U1290 ( .B(n1543), .A(n24), .Z(n27) );
  CNIVX2 U1291 ( .A(n1766), .Z(product[6]) );
  CNIVX1 U1292 ( .A(n1765), .Z(product[7]) );
  CANR1X2 U1293 ( .A(n204), .B(n1549), .C(n197), .Z(n195) );
  CIVX2 U1294 ( .A(n199), .Z(n197) );
  CEOX2 U1295 ( .A(a[14]), .B(n1745), .Z(n1393) );
  CENX4 U1296 ( .A(n1743), .B(a[14]), .Z(n66) );
  CENXL U1297 ( .A(n1710), .B(n1700), .Z(n1341) );
  CENXL U1298 ( .A(n1743), .B(n1700), .Z(n1173) );
  CENXL U1299 ( .A(n1727), .B(n1700), .Z(n1248) );
  CENXL U1300 ( .A(n1756), .B(n1700), .Z(n1101) );
  CENXL U1301 ( .A(n1754), .B(n1700), .Z(n1116) );
  CENXL U1302 ( .A(n1748), .B(n1700), .Z(n1133) );
  CENXL U1303 ( .A(n1525), .B(n1700), .Z(n1152) );
  CNIVX1 U1304 ( .A(n1378), .Z(n1696) );
  CIVXL U1305 ( .A(n221), .Z(n220) );
  CDLY1X2 U1306 ( .A(n1373), .Z(n1701) );
  CENXL U1307 ( .A(n1749), .B(n1369), .Z(n1128) );
  CENXL U1308 ( .A(n1737), .B(n1369), .Z(n1216) );
  CENXL U1309 ( .A(n1721), .B(n1369), .Z(n1272) );
  CENXL U1310 ( .A(n1716), .B(n1369), .Z(n1303) );
  CENXL U1311 ( .A(n1741), .B(n1369), .Z(n1191) );
  CENXL U1312 ( .A(n1745), .B(n1369), .Z(n1147) );
  CENXL U1313 ( .A(n1743), .B(n1369), .Z(n1168) );
  CENXL U1314 ( .A(n1728), .B(n1369), .Z(n1243) );
  CENXL U1315 ( .A(n1709), .B(n1361), .Z(n1328) );
  CENXL U1316 ( .A(n1735), .B(n1361), .Z(n1208) );
  CENXL U1317 ( .A(n1718), .B(n1361), .Z(n1264) );
  CENXL U1318 ( .A(n1712), .B(n1361), .Z(n1295) );
  CENXL U1319 ( .A(n1724), .B(n1361), .Z(n1235) );
  COND2XL U1320 ( .A(n77), .B(n1129), .C(n1128), .D(n74), .Z(n850) );
  COND2XL U1321 ( .A(n77), .B(n1752), .C(n1144), .D(n74), .Z(n785) );
  COND2XL U1322 ( .A(n77), .B(n1131), .C(n1130), .D(n74), .Z(n852) );
  COND2XL U1323 ( .A(n77), .B(n1130), .C(n1129), .D(n74), .Z(n851) );
  COND2XL U1324 ( .A(n77), .B(n1132), .C(n1131), .D(n74), .Z(n853) );
  COND2XL U1325 ( .A(n77), .B(n1142), .C(n1141), .D(n74), .Z(n863) );
  COND2XL U1326 ( .A(n77), .B(n1135), .C(n1134), .D(n74), .Z(n856) );
  COND2XL U1327 ( .A(n77), .B(n1133), .C(n1132), .D(n74), .Z(n854) );
  COND2XL U1328 ( .A(n77), .B(n1138), .C(n1137), .D(n74), .Z(n859) );
  COND2XL U1329 ( .A(n77), .B(n1137), .C(n74), .D(n1136), .Z(n858) );
  COND2XL U1330 ( .A(n77), .B(n1136), .C(n1135), .D(n74), .Z(n857) );
  COND2XL U1331 ( .A(n77), .B(n1134), .C(n1133), .D(n74), .Z(n855) );
  COND2XL U1332 ( .A(n77), .B(n1141), .C(n74), .D(n1140), .Z(n862) );
  COND2XL U1333 ( .A(n77), .B(n1139), .C(n74), .D(n1138), .Z(n860) );
  COND2XL U1334 ( .A(n77), .B(n1143), .C(n74), .D(n1142), .Z(n864) );
  COND2XL U1335 ( .A(n77), .B(n1140), .C(n1139), .D(n74), .Z(n861) );
  CANR1X1 U1336 ( .A(n260), .B(n268), .C(n261), .Z(n259) );
  CANR1XL U1337 ( .A(n208), .B(n180), .C(n181), .Z(n1533) );
  CANR1X2 U1338 ( .A(n190), .B(n1551), .C(n185), .Z(n183) );
  CENXL U1339 ( .A(n1746), .B(n1367), .Z(n1145) );
  CENXL U1340 ( .A(n1722), .B(n1367), .Z(n1270) );
  CENXL U1341 ( .A(n1711), .B(n1367), .Z(n1301) );
  CENXL U1342 ( .A(n1741), .B(n1367), .Z(n1189) );
  CENXL U1343 ( .A(n1737), .B(n1367), .Z(n1214) );
  CENXL U1344 ( .A(n1729), .B(n1367), .Z(n1241) );
  CIVX1 U1345 ( .A(n219), .Z(n217) );
  CNR2X1 U1346 ( .A(n182), .B(n194), .Z(n180) );
  COND1X1 U1347 ( .A(n195), .B(n182), .C(n183), .Z(n181) );
  CENXL U1348 ( .A(n1735), .B(n1365), .Z(n1212) );
  CENXL U1349 ( .A(n1718), .B(n1365), .Z(n1268) );
  CENXL U1350 ( .A(n1711), .B(n1365), .Z(n1299) );
  CENXL U1351 ( .A(n1709), .B(n1365), .Z(n1332) );
  CENXL U1352 ( .A(n1740), .B(n1365), .Z(n1187) );
  CENXL U1353 ( .A(n1724), .B(n1365), .Z(n1239) );
  CENXL U1354 ( .A(n158), .B(n121), .Z(product[29]) );
  COND1X1 U1355 ( .A(n209), .B(n221), .C(n210), .Z(n208) );
  COND1X1 U1356 ( .A(n259), .B(n242), .C(n243), .Z(n241) );
  CND2XL U1357 ( .A(n249), .B(n1558), .Z(n242) );
  CENX2 U1358 ( .A(n1740), .B(a[12]), .Z(n58) );
  CANR1XL U1359 ( .A(n1554), .B(n1537), .C(n155), .Z(n1534) );
  CANR1X1 U1360 ( .A(n1554), .B(n1537), .C(n155), .Z(n153) );
  COND2XL U1361 ( .A(n9), .B(n1347), .C(n6), .D(n1346), .Z(n1060) );
  CND2X4 U1362 ( .A(n1396), .B(n42), .Z(n44) );
  CIVX1 U1363 ( .A(n1731), .Z(n1727) );
  CENXL U1364 ( .A(n1542), .B(n150), .Z(product[31]) );
  CIVXL U1365 ( .A(n178), .Z(n1535) );
  CDLY1X2 U1366 ( .A(n1375), .Z(n1699) );
  CND2X1 U1367 ( .A(n1551), .B(n1546), .Z(n182) );
  CIVX2 U1368 ( .A(n21), .Z(n1723) );
  CENX2 U1369 ( .A(n1753), .B(a[20]), .Z(n89) );
  CIVX1 U1370 ( .A(n1755), .Z(n1753) );
  CND2X1 U1371 ( .A(n89), .B(n1390), .Z(n91) );
  CENXL U1372 ( .A(n1753), .B(n1693), .Z(n1124) );
  COND2X1 U1373 ( .A(n91), .B(n1110), .C(n1109), .D(n89), .Z(n833) );
  CND2X4 U1374 ( .A(n1400), .B(n6), .Z(n9) );
  CANR1XL U1375 ( .A(n1553), .B(n1540), .C(n163), .Z(n1536) );
  CENXL U1376 ( .A(n1527), .B(n1365), .Z(n1164) );
  CND2IXL U1377 ( .B(n1704), .A(n1527), .Z(n1184) );
  CENXL U1378 ( .A(n1703), .B(n1527), .Z(n1183) );
  CENXL U1379 ( .A(n1705), .B(n1527), .Z(n1182) );
  CENXL U1380 ( .A(n1695), .B(n1527), .Z(n1178) );
  CENXL U1381 ( .A(n1707), .B(n1527), .Z(n1180) );
  CENXL U1382 ( .A(n1527), .B(n1368), .Z(n1167) );
  CENXL U1383 ( .A(n1527), .B(n1367), .Z(n1166) );
  CENXL U1384 ( .A(n1527), .B(n1366), .Z(n1165) );
  COND2X1 U1385 ( .A(n69), .B(n1161), .C(n1160), .D(n66), .Z(n881) );
  CND2X4 U1386 ( .A(n1393), .B(n66), .Z(n69) );
  CDLY1X2 U1387 ( .A(n241), .Z(n1539) );
  COND1X1 U1388 ( .A(n167), .B(n179), .C(n168), .Z(n1540) );
  CIVXL U1389 ( .A(n1533), .Z(n178) );
  CIVX3 U1390 ( .A(n1528), .Z(n1710) );
  CENXL U1391 ( .A(n1710), .B(n1698), .Z(n1343) );
  CENXL U1392 ( .A(n1710), .B(n1695), .Z(n1346) );
  CENXL U1393 ( .A(n1710), .B(n1696), .Z(n1345) );
  CENXL U1394 ( .A(n1710), .B(n1369), .Z(n1336) );
  CENXL U1395 ( .A(n1710), .B(n1693), .Z(n1349) );
  CENXL U1396 ( .A(n1710), .B(n1704), .Z(n1351) );
  CENXL U1397 ( .A(n1710), .B(n1699), .Z(n1342) );
  COND2XL U1398 ( .A(n61), .B(n1165), .C(n1164), .D(n58), .Z(n884) );
  COND2XL U1399 ( .A(n61), .B(n1179), .C(n58), .D(n1178), .Z(n898) );
  COND2XL U1400 ( .A(n61), .B(n1169), .C(n1168), .D(n58), .Z(n888) );
  COND2XL U1401 ( .A(n61), .B(n1526), .C(n1184), .D(n58), .Z(n787) );
  COND2XL U1402 ( .A(n61), .B(n1172), .C(n1171), .D(n58), .Z(n891) );
  COND2XL U1403 ( .A(n61), .B(n1173), .C(n1172), .D(n58), .Z(n892) );
  COND2XL U1404 ( .A(n61), .B(n1183), .C(n58), .D(n1182), .Z(n902) );
  CNR2IXL U1405 ( .B(n1704), .A(n58), .Z(n903) );
  COND2XL U1406 ( .A(n61), .B(n1170), .C(n1169), .D(n58), .Z(n889) );
  COND2XL U1407 ( .A(n61), .B(n1171), .C(n1170), .D(n58), .Z(n890) );
  COND2XL U1408 ( .A(n61), .B(n1180), .C(n1179), .D(n58), .Z(n899) );
  COND2XL U1409 ( .A(n61), .B(n1182), .C(n1181), .D(n58), .Z(n901) );
  COND2XL U1410 ( .A(n61), .B(n1167), .C(n1166), .D(n58), .Z(n886) );
  COND2XL U1411 ( .A(n61), .B(n1168), .C(n1167), .D(n58), .Z(n887) );
  COND2XL U1412 ( .A(n61), .B(n1178), .C(n1177), .D(n58), .Z(n897) );
  COND2XL U1413 ( .A(n61), .B(n1177), .C(n1176), .D(n58), .Z(n896) );
  COND2XL U1414 ( .A(n61), .B(n1176), .C(n1175), .D(n58), .Z(n895) );
  COND2XL U1415 ( .A(n61), .B(n1175), .C(n1174), .D(n58), .Z(n894) );
  COND2XL U1416 ( .A(n61), .B(n1166), .C(n1165), .D(n58), .Z(n885) );
  COND2XL U1417 ( .A(n61), .B(n1174), .C(n1173), .D(n58), .Z(n893) );
  CND2IX2 U1418 ( .B(n1544), .A(n58), .Z(n61) );
  COND2XL U1419 ( .A(n36), .B(n1248), .C(n1247), .D(n33), .Z(n964) );
  COND2XL U1420 ( .A(n36), .B(n1251), .C(n1250), .D(n33), .Z(n967) );
  COND2XL U1421 ( .A(n36), .B(n1238), .C(n1237), .D(n33), .Z(n954) );
  COND2XL U1422 ( .A(n36), .B(n1234), .C(n1233), .D(n33), .Z(n950) );
  COND2XL U1423 ( .A(n36), .B(n1246), .C(n1245), .D(n33), .Z(n962) );
  COND2XL U1424 ( .A(n36), .B(n1254), .C(n1253), .D(n33), .Z(n970) );
  COND2XL U1425 ( .A(n36), .B(n1247), .C(n1246), .D(n33), .Z(n963) );
  COND2XL U1426 ( .A(n36), .B(n1252), .C(n1251), .D(n33), .Z(n968) );
  COND2XL U1427 ( .A(n36), .B(n1237), .C(n1236), .D(n33), .Z(n953) );
  COND2XL U1428 ( .A(n36), .B(n1242), .C(n1241), .D(n33), .Z(n958) );
  COND2XL U1429 ( .A(n36), .B(n1241), .C(n1240), .D(n33), .Z(n957) );
  COND2XL U1430 ( .A(n36), .B(n1236), .C(n1235), .D(n33), .Z(n952) );
  COND2XL U1431 ( .A(n36), .B(n1255), .C(n1254), .D(n33), .Z(n971) );
  COND2XL U1432 ( .A(n36), .B(n1243), .C(n1242), .D(n33), .Z(n959) );
  COND2XL U1433 ( .A(n36), .B(n1235), .C(n1234), .D(n33), .Z(n951) );
  COND2XL U1434 ( .A(n36), .B(n1249), .C(n1248), .D(n33), .Z(n965) );
  COND2XL U1435 ( .A(n36), .B(n1245), .C(n1244), .D(n33), .Z(n961) );
  COND2XL U1436 ( .A(n36), .B(n1244), .C(n1243), .D(n33), .Z(n960) );
  COND2XL U1437 ( .A(n36), .B(n1240), .C(n1239), .D(n33), .Z(n956) );
  COND2XL U1438 ( .A(n36), .B(n1239), .C(n1238), .D(n33), .Z(n955) );
  COND2XL U1439 ( .A(n36), .B(n1256), .C(n33), .D(n1255), .Z(n972) );
  COND2XL U1440 ( .A(n36), .B(n1253), .C(n1252), .D(n33), .Z(n969) );
  COND2XL U1441 ( .A(n36), .B(n1258), .C(n33), .D(n1257), .Z(n974) );
  CENXL U1442 ( .A(n1720), .B(n1372), .Z(n1275) );
  CENXL U1443 ( .A(n1720), .B(n1698), .Z(n1279) );
  COND2XL U1444 ( .A(n36), .B(n1257), .C(n1256), .D(n33), .Z(n973) );
  COND2XL U1445 ( .A(n36), .B(n1730), .C(n1259), .D(n33), .Z(n790) );
  CENXL U1446 ( .A(n1720), .B(n1701), .Z(n1276) );
  COND1X1 U1447 ( .A(n151), .B(n153), .C(n152), .Z(n150) );
  CNIVX1 U1448 ( .A(n1381), .Z(n1707) );
  CNIVX1 U1449 ( .A(n1377), .Z(n1697) );
  CENXL U1450 ( .A(n1529), .B(n1702), .Z(n1338) );
  CND2IXL U1451 ( .B(n1704), .A(n1529), .Z(n1352) );
  CENXL U1452 ( .A(n1529), .B(n1366), .Z(n1333) );
  CENXL U1453 ( .A(n1529), .B(n1367), .Z(n1334) );
  CENXL U1454 ( .A(n1529), .B(n1368), .Z(n1335) );
  CENXL U1455 ( .A(n1705), .B(n1529), .Z(n1350) );
  CENXL U1456 ( .A(n1707), .B(n1529), .Z(n1348) );
  CENXL U1457 ( .A(n1529), .B(n1370), .Z(n1337) );
  CENXL U1458 ( .A(n1710), .B(n1694), .Z(n1347) );
  CENXL U1459 ( .A(n1694), .B(n1763), .Z(n1083) );
  CENXL U1460 ( .A(n1747), .B(n1694), .Z(n1139) );
  COND1X1 U1461 ( .A(n159), .B(n161), .C(n160), .Z(n1537) );
  COAN1XL U1462 ( .A(n209), .B(n221), .C(n210), .Z(n1538) );
  CANR1X1 U1463 ( .A(n1553), .B(n1540), .C(n163), .Z(n161) );
  CNR2XL U1464 ( .A(n251), .B(n256), .Z(n249) );
  CIVX1 U1465 ( .A(n1528), .Z(n1709) );
  COND2XL U1466 ( .A(n97), .B(n1091), .C(n1090), .D(n95), .Z(n815) );
  CIVX1 U1467 ( .A(a[0]), .Z(n6) );
  COR2XL U1468 ( .A(n1567), .B(n1565), .Z(n1560) );
  CANR1XL U1469 ( .A(n1691), .B(n286), .C(n283), .Z(n281) );
  CANR1XL U1470 ( .A(n1685), .B(n1690), .C(n291), .Z(n289) );
  CNR2XL U1471 ( .A(n224), .B(n227), .Z(n222) );
  CANR1XL U1472 ( .A(n302), .B(n1556), .C(n299), .Z(n297) );
  CND2XL U1473 ( .A(n340), .B(n304), .Z(n147) );
  CENX1 U1474 ( .A(n1709), .B(n1697), .Z(n1344) );
  CIVX2 U1475 ( .A(n1762), .Z(n1761) );
  COND2X1 U1476 ( .A(n1095), .B(n97), .C(n1094), .D(n95), .Z(n819) );
  CNR2IX1 U1477 ( .B(n1704), .A(n42), .Z(n949) );
  COND2X1 U1478 ( .A(n53), .B(n1203), .C(n1202), .D(n50), .Z(n921) );
  COND2X1 U1479 ( .A(n1080), .B(n100), .C(n1081), .D(n102), .Z(n806) );
  CENXL U1480 ( .A(a[12]), .B(n1527), .Z(n1544) );
  CNIVX1 U1481 ( .A(n1382), .Z(n1693) );
  CNIVX1 U1482 ( .A(n1376), .Z(n1698) );
  CND2X1 U1483 ( .A(n95), .B(n1389), .Z(n97) );
  CEOXL U1484 ( .A(a[18]), .B(n1754), .Z(n1391) );
  CIVX1 U1485 ( .A(n113), .Z(n1410) );
  CANR1X1 U1486 ( .A(n208), .B(n180), .C(n181), .Z(n179) );
  CND2XL U1487 ( .A(n1550), .B(n1547), .Z(n209) );
  CEOXL U1488 ( .A(n1534), .B(n120), .Z(product[30]) );
  CEOXL U1489 ( .A(n124), .B(n173), .Z(product[26]) );
  CND2XL U1490 ( .A(n1552), .B(n172), .Z(n124) );
  CEOXL U1491 ( .A(n126), .B(n188), .Z(product[24]) );
  CND2XL U1492 ( .A(n1551), .B(n187), .Z(n126) );
  CEOXL U1493 ( .A(n130), .B(n215), .Z(product[20]) );
  CND2XL U1494 ( .A(n1550), .B(n214), .Z(n130) );
  CND2XL U1495 ( .A(n315), .B(n160), .Z(n122) );
  CND2XL U1496 ( .A(n322), .B(n202), .Z(n129) );
  CEOXL U1497 ( .A(n297), .B(n145), .Z(product[5]) );
  CEOXL U1498 ( .A(n305), .B(n147), .Z(product[3]) );
  CND2XL U1499 ( .A(n1556), .B(n301), .Z(n146) );
  CND2XL U1500 ( .A(n1555), .B(n309), .Z(n148) );
  CND2XL U1501 ( .A(n1554), .B(n157), .Z(n121) );
  CND2XL U1502 ( .A(n1553), .B(n165), .Z(n123) );
  CND2XL U1503 ( .A(n1548), .B(n177), .Z(n125) );
  CND2XL U1504 ( .A(n1546), .B(n192), .Z(n127) );
  CND2XL U1505 ( .A(n1547), .B(n219), .Z(n131) );
  CND2XL U1506 ( .A(n1549), .B(n322), .Z(n194) );
  CND2XL U1507 ( .A(n755), .B(n760), .Z(n285) );
  CNR2XL U1508 ( .A(n262), .B(n265), .Z(n260) );
  CND2XL U1509 ( .A(n332), .B(n266), .Z(n139) );
  CND2XL U1510 ( .A(n1558), .B(n247), .Z(n135) );
  CND2XL U1511 ( .A(n327), .B(n235), .Z(n134) );
  CND2XL U1512 ( .A(n330), .B(n257), .Z(n137) );
  CND2XL U1513 ( .A(n1559), .B(n232), .Z(n133) );
  CND2XL U1514 ( .A(n325), .B(n225), .Z(n132) );
  CND2XL U1515 ( .A(n777), .B(n792), .Z(n304) );
  CND2XL U1516 ( .A(n1559), .B(n327), .Z(n227) );
  CNR2XL U1517 ( .A(n761), .B(n766), .Z(n287) );
  COR2XL U1518 ( .A(n1063), .B(n1033), .Z(n1555) );
  CND2XL U1519 ( .A(n767), .B(n770), .Z(n293) );
  COR2XL U1520 ( .A(n1064), .B(n793), .Z(n1541) );
  CENX1 U1521 ( .A(n343), .B(n358), .Z(n1542) );
  CND2XL U1522 ( .A(n695), .B(n706), .Z(n252) );
  CND2XL U1523 ( .A(n1561), .B(n274), .Z(n140) );
  CNR2IXL U1524 ( .B(n1704), .A(n74), .Z(n865) );
  CNR2IXL U1525 ( .B(n1704), .A(n95), .Z(n823) );
  CNR2IXL U1526 ( .B(n1704), .A(n105), .Z(n805) );
  CND2XL U1527 ( .A(n1560), .B(n279), .Z(n141) );
  CNR2IXL U1528 ( .B(n1704), .A(n33), .Z(n975) );
  COND2XL U1529 ( .A(n18), .B(n1315), .C(n15), .D(n1314), .Z(n1029) );
  CNR2IXL U1530 ( .B(n1704), .A(n100), .Z(n813) );
  COND2XL U1531 ( .A(n1097), .B(n97), .C(n1096), .D(n95), .Z(n821) );
  CNR2IXL U1532 ( .B(n1704), .A(n110), .Z(n799) );
  COND2XL U1533 ( .A(n1093), .B(n97), .C(n1092), .D(n95), .Z(n817) );
  CNR2IXL U1534 ( .B(n1704), .A(n66), .Z(n883) );
  CND2XL U1535 ( .A(n719), .B(n728), .Z(n263) );
  CEOXL U1536 ( .A(n778), .B(n806), .Z(n357) );
  CNR2IXL U1537 ( .B(n1704), .A(n6), .Z(product[0]) );
  CNIVXL U1538 ( .A(n1374), .Z(n1700) );
  CENXL U1539 ( .A(a[4]), .B(n1722), .Z(n1543) );
  CIVX3 U1540 ( .A(n1564), .Z(n42) );
  CIVX3 U1541 ( .A(n1562), .Z(n24) );
  CEOXL U1542 ( .A(a[16]), .B(n1749), .Z(n1392) );
  CNIVXL U1543 ( .A(n1381), .Z(n1708) );
  CND2IXL U1544 ( .B(n1704), .A(n109), .Z(n1072) );
  CND2IXL U1545 ( .B(n1704), .A(n113), .Z(n1067) );
  COND1XL U1546 ( .A(n194), .B(n1538), .C(n195), .Z(n193) );
  CANR1XL U1547 ( .A(n310), .B(n1555), .C(n307), .Z(n305) );
  CND2X1 U1548 ( .A(n1552), .B(n1548), .Z(n167) );
  COND1XL U1549 ( .A(n159), .B(n1536), .C(n160), .Z(n158) );
  COND1XL U1550 ( .A(n305), .B(n303), .C(n304), .Z(n302) );
  CANR1XL U1551 ( .A(n1547), .B(n220), .C(n217), .Z(n215) );
  CENX1 U1552 ( .A(n200), .B(n128), .Z(product[22]) );
  CND2X1 U1553 ( .A(n1549), .B(n199), .Z(n128) );
  COND1XL U1554 ( .A(n201), .B(n1538), .C(n202), .Z(n200) );
  CENX1 U1555 ( .A(n146), .B(n302), .Z(product[4]) );
  CENX1 U1556 ( .A(n193), .B(n127), .Z(product[23]) );
  CENX1 U1557 ( .A(n178), .B(n125), .Z(product[25]) );
  CENX1 U1558 ( .A(n166), .B(n123), .Z(product[27]) );
  CENX1 U1559 ( .A(n220), .B(n131), .Z(product[19]) );
  COND1XL U1560 ( .A(n297), .B(n295), .C(n296), .Z(n294) );
  CND2X1 U1561 ( .A(n338), .B(n296), .Z(n145) );
  CND2X1 U1562 ( .A(n313), .B(n152), .Z(n120) );
  CEOXL U1563 ( .A(n122), .B(n1536), .Z(product[28]) );
  CANR1XL U1564 ( .A(n1548), .B(n178), .C(n175), .Z(n173) );
  CANR1XL U1565 ( .A(n1546), .B(n193), .C(n190), .Z(n188) );
  CEOXL U1566 ( .A(n129), .B(n1538), .Z(product[21]) );
  CENX1 U1567 ( .A(n148), .B(n310), .Z(product[2]) );
  COR2X1 U1568 ( .A(n755), .B(n760), .Z(n1545) );
  CEOX1 U1569 ( .A(n135), .B(n248), .Z(product[15]) );
  CANR1XL U1570 ( .A(n249), .B(n258), .C(n250), .Z(n248) );
  COND1XL U1571 ( .A(n266), .B(n262), .C(n263), .Z(n261) );
  COND1XL U1572 ( .A(n228), .B(n224), .C(n225), .Z(n223) );
  CENX1 U1573 ( .A(n264), .B(n138), .Z(product[12]) );
  CND2X1 U1574 ( .A(n331), .B(n263), .Z(n138) );
  COND1XL U1575 ( .A(n265), .B(n267), .C(n266), .Z(n264) );
  CENX1 U1576 ( .A(n258), .B(n137), .Z(product[13]) );
  CENX1 U1577 ( .A(n233), .B(n133), .Z(product[17]) );
  COND1XL U1578 ( .A(n234), .B(n240), .C(n235), .Z(n233) );
  CENX1 U1579 ( .A(n226), .B(n132), .Z(product[18]) );
  COND1XL U1580 ( .A(n227), .B(n240), .C(n228), .Z(n226) );
  CNR2X1 U1581 ( .A(n579), .B(n598), .Z(n201) );
  CNR2X1 U1582 ( .A(n415), .B(n440), .Z(n159) );
  CNR2X1 U1583 ( .A(n359), .B(n386), .Z(n151) );
  CNR2X1 U1584 ( .A(n771), .B(n774), .Z(n295) );
  CNR2X1 U1585 ( .A(n777), .B(n792), .Z(n303) );
  CEOX1 U1586 ( .A(n139), .B(n267), .Z(product[11]) );
  CEOX1 U1587 ( .A(n136), .B(n253), .Z(product[14]) );
  CND2X1 U1588 ( .A(n329), .B(n252), .Z(n136) );
  CANR1XL U1589 ( .A(n330), .B(n258), .C(n255), .Z(n253) );
  CEOX1 U1590 ( .A(n134), .B(n240), .Z(product[16]) );
  COR2X1 U1591 ( .A(n537), .B(n558), .Z(n1546) );
  COR2X1 U1592 ( .A(n617), .B(n634), .Z(n1547) );
  COR2X1 U1593 ( .A(n491), .B(n514), .Z(n1548) );
  COR2X1 U1594 ( .A(n559), .B(n578), .Z(n1549) );
  COR2X1 U1595 ( .A(n599), .B(n616), .Z(n1550) );
  CND2X1 U1596 ( .A(n579), .B(n598), .Z(n202) );
  COR2X1 U1597 ( .A(n515), .B(n536), .Z(n1551) );
  COR2X1 U1598 ( .A(n467), .B(n490), .Z(n1552) );
  CND2X1 U1599 ( .A(n537), .B(n558), .Z(n192) );
  CND2X1 U1600 ( .A(n617), .B(n634), .Z(n219) );
  CND2X1 U1601 ( .A(n515), .B(n536), .Z(n187) );
  CND2X1 U1602 ( .A(n559), .B(n578), .Z(n199) );
  CND2X1 U1603 ( .A(n599), .B(n616), .Z(n214) );
  CND2X1 U1604 ( .A(n491), .B(n514), .Z(n177) );
  CND2X1 U1605 ( .A(n1064), .B(n793), .Z(n312) );
  CND2X1 U1606 ( .A(n467), .B(n490), .Z(n172) );
  CND2X1 U1607 ( .A(n441), .B(n466), .Z(n165) );
  CND2X1 U1608 ( .A(n1063), .B(n1033), .Z(n309) );
  CND2X1 U1609 ( .A(n775), .B(n776), .Z(n301) );
  CND2X1 U1610 ( .A(n387), .B(n414), .Z(n157) );
  CND2X1 U1611 ( .A(n771), .B(n774), .Z(n296) );
  CND2X1 U1612 ( .A(n415), .B(n440), .Z(n160) );
  CND2X1 U1613 ( .A(n359), .B(n386), .Z(n152) );
  COR2X1 U1614 ( .A(n441), .B(n466), .Z(n1553) );
  COR2X1 U1615 ( .A(n387), .B(n414), .Z(n1554) );
  COR2X1 U1616 ( .A(n775), .B(n776), .Z(n1556) );
  CND2XL U1617 ( .A(n761), .B(n766), .Z(n288) );
  COR2X1 U1618 ( .A(n767), .B(n770), .Z(n1557) );
  CIVX2 U1619 ( .A(n1764), .Z(n1763) );
  CENX1 U1620 ( .A(n1701), .B(n1757), .Z(n1100) );
  CENX1 U1621 ( .A(n1702), .B(n1523), .Z(n1113) );
  COND1XL U1622 ( .A(n281), .B(n269), .C(n270), .Z(n268) );
  CND2X1 U1623 ( .A(n1561), .B(n1560), .Z(n269) );
  CANR1XL U1624 ( .A(n277), .B(n1561), .C(n272), .Z(n270) );
  CIVX2 U1625 ( .A(n1526), .Z(n1743) );
  CIVX2 U1626 ( .A(n1742), .Z(n1740) );
  CENX1 U1627 ( .A(n1699), .B(n1761), .Z(n1089) );
  CNR2X1 U1628 ( .A(n729), .B(n738), .Z(n265) );
  CNR2X1 U1629 ( .A(n695), .B(n706), .Z(n251) );
  CNR2X1 U1630 ( .A(n635), .B(n650), .Z(n224) );
  CNR2X1 U1631 ( .A(n719), .B(n728), .Z(n262) );
  CNR2IXL U1632 ( .B(n1704), .A(n15), .Z(n1033) );
  CENX1 U1633 ( .A(n1761), .B(n1693), .Z(n1096) );
  CENX1 U1634 ( .A(n1761), .B(n1694), .Z(n1094) );
  CENX1 U1635 ( .A(n1693), .B(n1763), .Z(n1085) );
  CENX1 U1636 ( .A(n1696), .B(n1763), .Z(n1081) );
  CENX1 U1637 ( .A(n1734), .B(n1698), .Z(n1223) );
  CENX1 U1638 ( .A(n1744), .B(n1693), .Z(n1160) );
  CENX1 U1639 ( .A(n1744), .B(n1694), .Z(n1158) );
  CENX1 U1640 ( .A(n1747), .B(n1693), .Z(n1141) );
  CENX1 U1641 ( .A(n1744), .B(n1696), .Z(n1156) );
  CENX1 U1642 ( .A(n1743), .B(n1699), .Z(n1174) );
  CENX1 U1643 ( .A(n1697), .B(n1746), .Z(n1155) );
  CENX1 U1644 ( .A(n1747), .B(n1696), .Z(n1137) );
  CENX1 U1645 ( .A(n1754), .B(n1694), .Z(n1122) );
  CENX1 U1646 ( .A(n1757), .B(n1693), .Z(n1109) );
  CENX1 U1647 ( .A(n1744), .B(n1698), .Z(n1154) );
  CENX1 U1648 ( .A(n1525), .B(n1699), .Z(n1153) );
  CENX1 U1649 ( .A(n1747), .B(n1698), .Z(n1135) );
  CENX1 U1650 ( .A(n1757), .B(n1694), .Z(n1107) );
  CENX1 U1651 ( .A(n1699), .B(n1750), .Z(n1134) );
  CENX1 U1652 ( .A(n1525), .B(n1701), .Z(n1151) );
  CENX1 U1653 ( .A(n1756), .B(n1696), .Z(n1105) );
  CENX1 U1654 ( .A(n1756), .B(n1698), .Z(n1103) );
  CENX1 U1655 ( .A(n1701), .B(n1523), .Z(n1115) );
  CENX1 U1656 ( .A(n1726), .B(n1695), .Z(n1253) );
  CENX1 U1657 ( .A(n1726), .B(n1694), .Z(n1254) );
  CENX1 U1658 ( .A(n1733), .B(n1693), .Z(n1229) );
  CENX1 U1659 ( .A(n1733), .B(n1694), .Z(n1227) );
  CENX1 U1660 ( .A(n1725), .B(n1696), .Z(n1252) );
  CENX1 U1661 ( .A(n1728), .B(n1698), .Z(n1250) );
  CENX1 U1662 ( .A(n1740), .B(n1699), .Z(n1197) );
  CENX1 U1663 ( .A(n1754), .B(n1698), .Z(n1118) );
  CENX1 U1664 ( .A(n1726), .B(n1693), .Z(n1256) );
  CENX1 U1665 ( .A(n1733), .B(n1697), .Z(n1224) );
  CENX1 U1666 ( .A(n1733), .B(n1696), .Z(n1225) );
  CENX1 U1667 ( .A(n1728), .B(n1699), .Z(n1249) );
  CENX1 U1668 ( .A(n1740), .B(n1694), .Z(n1202) );
  CENX1 U1669 ( .A(n1743), .B(n1693), .Z(n1181) );
  CENX1 U1670 ( .A(n1740), .B(n1696), .Z(n1200) );
  CENX1 U1671 ( .A(n1735), .B(n1699), .Z(n1222) );
  CENX1 U1672 ( .A(n1743), .B(n1696), .Z(n1177) );
  CENX1 U1673 ( .A(n1743), .B(n1697), .Z(n1176) );
  CENX1 U1674 ( .A(n1743), .B(n1698), .Z(n1175) );
  CENX1 U1675 ( .A(n1740), .B(n1701), .Z(n1195) );
  CENX1 U1676 ( .A(n1743), .B(n1702), .Z(n1170) );
  CENX1 U1677 ( .A(n1748), .B(n1701), .Z(n1132) );
  CENX1 U1678 ( .A(n1745), .B(n1702), .Z(n1149) );
  CENX1 U1679 ( .A(n1761), .B(n1696), .Z(n1092) );
  CENX1 U1680 ( .A(n1749), .B(n1702), .Z(n1130) );
  CENX1 U1681 ( .A(n1761), .B(n1698), .Z(n1090) );
  CENX1 U1682 ( .A(n1740), .B(n1693), .Z(n1204) );
  CENX1 U1683 ( .A(n1695), .B(n1733), .Z(n1226) );
  CENX1 U1684 ( .A(n1725), .B(n1697), .Z(n1251) );
  CENX1 U1685 ( .A(n1743), .B(n1694), .Z(n1179) );
  CENX1 U1686 ( .A(n1740), .B(n1697), .Z(n1199) );
  CENX1 U1687 ( .A(n1724), .B(n1701), .Z(n1247) );
  CENX1 U1688 ( .A(n1740), .B(n1698), .Z(n1198) );
  CENX1 U1689 ( .A(n1728), .B(n1702), .Z(n1245) );
  CENX1 U1690 ( .A(n1736), .B(n1701), .Z(n1220) );
  CENX1 U1691 ( .A(n1736), .B(n1702), .Z(n1218) );
  CENX1 U1692 ( .A(n1741), .B(n1702), .Z(n1193) );
  CENX1 U1693 ( .A(n1743), .B(n1701), .Z(n1172) );
  CENX1 U1694 ( .A(n1705), .B(n1715), .Z(n1317) );
  CENX1 U1695 ( .A(n1716), .B(n1696), .Z(n1312) );
  CENX1 U1696 ( .A(n1719), .B(n1697), .Z(n1280) );
  CENX1 U1697 ( .A(n1715), .B(n1699), .Z(n1309) );
  CENX1 U1698 ( .A(n1705), .B(n1746), .Z(n1161) );
  CENX1 U1699 ( .A(n1705), .B(n1750), .Z(n1142) );
  CENX1 U1700 ( .A(n1707), .B(n1746), .Z(n1159) );
  CENX1 U1701 ( .A(n1707), .B(n1750), .Z(n1140) );
  CENX1 U1702 ( .A(n1705), .B(n1523), .Z(n1125) );
  CENX1 U1703 ( .A(n1695), .B(n1746), .Z(n1157) );
  CENX1 U1704 ( .A(n1705), .B(n1758), .Z(n1110) );
  CENX1 U1705 ( .A(n1707), .B(n1523), .Z(n1123) );
  CENX1 U1706 ( .A(n1695), .B(n1523), .Z(n1121) );
  CENX1 U1707 ( .A(n1707), .B(n1758), .Z(n1108) );
  CENX1 U1708 ( .A(n1695), .B(n1758), .Z(n1106) );
  CENX1 U1709 ( .A(n1697), .B(n1523), .Z(n1119) );
  CENX1 U1710 ( .A(n1697), .B(n1758), .Z(n1104) );
  CENX1 U1711 ( .A(n1699), .B(n1758), .Z(n1102) );
  CENX1 U1712 ( .A(n1707), .B(n1716), .Z(n1315) );
  CENX1 U1713 ( .A(n1719), .B(n1693), .Z(n1285) );
  CENX1 U1714 ( .A(n1718), .B(n1695), .Z(n1282) );
  CENX1 U1715 ( .A(n1719), .B(n1696), .Z(n1281) );
  CENX1 U1716 ( .A(n1715), .B(n1697), .Z(n1311) );
  CENX1 U1717 ( .A(n1714), .B(n1698), .Z(n1310) );
  CENX1 U1718 ( .A(n1719), .B(n1699), .Z(n1278) );
  CENX1 U1719 ( .A(n1714), .B(n1701), .Z(n1307) );
  CENX1 U1720 ( .A(n1699), .B(n1523), .Z(n1117) );
  CENX1 U1721 ( .A(n1713), .B(n1694), .Z(n1314) );
  CENX1 U1722 ( .A(n1713), .B(n1695), .Z(n1313) );
  CENX1 U1723 ( .A(n1713), .B(n1693), .Z(n1316) );
  CENX1 U1724 ( .A(n1705), .B(n1729), .Z(n1257) );
  CENX1 U1725 ( .A(n1707), .B(n1721), .Z(n1284) );
  CENX1 U1726 ( .A(n1705), .B(n1737), .Z(n1230) );
  CENX1 U1727 ( .A(n1710), .B(n1701), .Z(n1340) );
  CENX1 U1728 ( .A(n1716), .B(n1702), .Z(n1305) );
  CENX1 U1729 ( .A(n1721), .B(n1702), .Z(n1274) );
  CENX1 U1730 ( .A(n1695), .B(n1751), .Z(n1138) );
  CENX1 U1731 ( .A(n1697), .B(n1751), .Z(n1136) );
  CENX1 U1732 ( .A(n1697), .B(n1761), .Z(n1091) );
  CENX1 U1733 ( .A(n1705), .B(n1718), .Z(n1286) );
  CENX1 U1734 ( .A(n1707), .B(n1729), .Z(n1255) );
  CENX1 U1735 ( .A(n1707), .B(n1735), .Z(n1228) );
  CENX1 U1736 ( .A(n1707), .B(n1741), .Z(n1203) );
  CENX1 U1737 ( .A(n1705), .B(n1761), .Z(n1097) );
  CENX1 U1738 ( .A(n1707), .B(n1761), .Z(n1095) );
  CENX1 U1739 ( .A(n1705), .B(n1763), .Z(n1086) );
  CENX1 U1740 ( .A(n1695), .B(n1761), .Z(n1093) );
  CENX1 U1741 ( .A(n1707), .B(n1763), .Z(n1084) );
  CENX1 U1742 ( .A(n1695), .B(n1763), .Z(n1082) );
  CNR2X1 U1743 ( .A(n707), .B(n718), .Z(n256) );
  CENX1 U1744 ( .A(n1703), .B(n1761), .Z(n1098) );
  CENX1 U1745 ( .A(n1726), .B(n1704), .Z(n1258) );
  CENX1 U1746 ( .A(n1734), .B(n1703), .Z(n1231) );
  CENX1 U1747 ( .A(n1703), .B(n1746), .Z(n1162) );
  CENX1 U1748 ( .A(n1703), .B(n1750), .Z(n1143) );
  CENX1 U1749 ( .A(n1703), .B(n1523), .Z(n1126) );
  CENX1 U1750 ( .A(n1703), .B(n1741), .Z(n1206) );
  CENX1 U1751 ( .A(n1703), .B(n1758), .Z(n1111) );
  CENX1 U1752 ( .A(n1703), .B(n1763), .Z(n1087) );
  CENX1 U1753 ( .A(n1697), .B(n1763), .Z(n1080) );
  CENX1 U1754 ( .A(n1719), .B(n1704), .Z(n1287) );
  CNR2IX1 U1755 ( .B(n1704), .A(n24), .Z(n1003) );
  CENX1 U1756 ( .A(n1714), .B(n1703), .Z(n1318) );
  CNR2X1 U1757 ( .A(n667), .B(n680), .Z(n234) );
  CNR2IX1 U1758 ( .B(n1704), .A(n114), .Z(n795) );
  CEOX1 U1759 ( .A(n275), .B(n140), .Z(product[10]) );
  CANR1XL U1760 ( .A(n1560), .B(n280), .C(n277), .Z(n275) );
  CNR2IX1 U1761 ( .B(n1704), .A(n82), .Z(n849) );
  COR2X1 U1762 ( .A(n681), .B(n694), .Z(n1558) );
  COR2X1 U1763 ( .A(n651), .B(n666), .Z(n1559) );
  CND2X1 U1764 ( .A(n667), .B(n680), .Z(n235) );
  CNR2IX1 U1765 ( .B(n1704), .A(n89), .Z(n835) );
  CND2X1 U1766 ( .A(n707), .B(n718), .Z(n257) );
  CNR2IXL U1767 ( .B(n1704), .A(n50), .Z(n925) );
  CND2X1 U1768 ( .A(n729), .B(n738), .Z(n266) );
  CND2X1 U1769 ( .A(n651), .B(n666), .Z(n232) );
  CND2X1 U1770 ( .A(n681), .B(n694), .Z(n247) );
  CND2X1 U1771 ( .A(n635), .B(n650), .Z(n225) );
  CENX1 U1772 ( .A(n141), .B(n280), .Z(product[9]) );
  CENX1 U1773 ( .A(n1525), .B(a[16]), .Z(n74) );
  CENX1 U1774 ( .A(n1756), .B(a[22]), .Z(n95) );
  CENX1 U1775 ( .A(n1761), .B(a[24]), .Z(n100) );
  CENX1 U1776 ( .A(n1763), .B(a[26]), .Z(n105) );
  CENX1 U1777 ( .A(n1748), .B(n1372), .Z(n1131) );
  CENX1 U1778 ( .A(n1753), .B(n1372), .Z(n1114) );
  CENX1 U1779 ( .A(n1745), .B(n1372), .Z(n1150) );
  CENX1 U1780 ( .A(n1727), .B(n1372), .Z(n1246) );
  CENX1 U1781 ( .A(n1736), .B(n1372), .Z(n1219) );
  CENX1 U1782 ( .A(n1743), .B(n1372), .Z(n1171) );
  CENX1 U1783 ( .A(n1725), .B(n1363), .Z(n1237) );
  CENX1 U1784 ( .A(n1736), .B(n1363), .Z(n1210) );
  CENX1 U1785 ( .A(n1711), .B(n1363), .Z(n1297) );
  CENX1 U1786 ( .A(n1715), .B(n1372), .Z(n1306) );
  CENX1 U1787 ( .A(n1722), .B(n1368), .Z(n1271) );
  CENX1 U1788 ( .A(n1709), .B(n1363), .Z(n1330) );
  CENX1 U1789 ( .A(n1718), .B(n1363), .Z(n1266) );
  CENX1 U1790 ( .A(n1710), .B(n1372), .Z(n1339) );
  CENX1 U1791 ( .A(n104), .B(a[28]), .Z(n110) );
  COND1XL U1792 ( .A(n1688), .B(n289), .C(n1687), .Z(n286) );
  CENX1 U1793 ( .A(n1727), .B(b[25]), .Z(n1233) );
  CENX1 U1794 ( .A(n1719), .B(b[27]), .Z(n1260) );
  CENX1 U1795 ( .A(n1708), .B(n109), .Z(n1068) );
  CENX1 U1796 ( .A(n109), .B(a[30]), .Z(n114) );
  CENX1 U1797 ( .A(n1713), .B(b[29]), .Z(n1289) );
  CNIVX1 U1798 ( .A(n1383), .Z(n1705) );
  CEOX1 U1799 ( .A(a[0]), .B(n1529), .Z(n1400) );
  CND2X2 U1800 ( .A(n1397), .B(n33), .Z(n36) );
  CEOX1 U1801 ( .A(a[6]), .B(n1729), .Z(n1397) );
  CENX1 U1802 ( .A(n1740), .B(n1363), .Z(n1185) );
  CENX1 U1803 ( .A(n1695), .B(n104), .Z(n1073) );
  CENX1 U1804 ( .A(n1703), .B(n113), .Z(n1066) );
  CENX1 U1805 ( .A(n1706), .B(n113), .Z(n1065) );
  CEOX1 U1806 ( .A(a[8]), .B(n1737), .Z(n1396) );
  CENX1 U1807 ( .A(n1728), .B(n1370), .Z(n1244) );
  CENX1 U1808 ( .A(n1735), .B(n1370), .Z(n1217) );
  CENX1 U1809 ( .A(n1734), .B(n1364), .Z(n1211) );
  CENX1 U1810 ( .A(n1745), .B(n1370), .Z(n1148) );
  CENX1 U1811 ( .A(n1749), .B(n1370), .Z(n1129) );
  CENX1 U1812 ( .A(n1740), .B(n1364), .Z(n1186) );
  CENX1 U1813 ( .A(n1735), .B(n1362), .Z(n1209) );
  CENX1 U1814 ( .A(n1724), .B(b[24]), .Z(n1234) );
  CENX1 U1815 ( .A(n1743), .B(n1370), .Z(n1169) );
  CENX1 U1816 ( .A(n1725), .B(n1364), .Z(n1238) );
  CENX1 U1817 ( .A(n1724), .B(n1362), .Z(n1236) );
  CENX1 U1818 ( .A(n1693), .B(n104), .Z(n1076) );
  CENX1 U1819 ( .A(n1693), .B(n109), .Z(n1069) );
  CENX1 U1820 ( .A(n1711), .B(b[26]), .Z(n1292) );
  CENX1 U1821 ( .A(n1718), .B(b[25]), .Z(n1262) );
  CENX1 U1822 ( .A(n1711), .B(b[27]), .Z(n1291) );
  CENX1 U1823 ( .A(n1719), .B(b[26]), .Z(n1261) );
  CENX1 U1824 ( .A(n1711), .B(b[28]), .Z(n1290) );
  CENX1 U1825 ( .A(n1716), .B(n1370), .Z(n1304) );
  CENX1 U1826 ( .A(n1722), .B(n1370), .Z(n1273) );
  CENX1 U1827 ( .A(n1709), .B(n1364), .Z(n1331) );
  CENX1 U1828 ( .A(n1711), .B(n1364), .Z(n1298) );
  CENX1 U1829 ( .A(n1712), .B(n1362), .Z(n1296) );
  CENX1 U1830 ( .A(n1718), .B(n1364), .Z(n1267) );
  CENX1 U1831 ( .A(n1709), .B(b[25]), .Z(n1326) );
  CENX1 U1832 ( .A(n1718), .B(n1362), .Z(n1265) );
  CENX1 U1833 ( .A(n1718), .B(b[24]), .Z(n1263) );
  CENX1 U1834 ( .A(n1709), .B(b[28]), .Z(n1323) );
  CENX1 U1835 ( .A(n1709), .B(b[29]), .Z(n1322) );
  CENX1 U1836 ( .A(n1709), .B(b[30]), .Z(n1321) );
  CENX1 U1837 ( .A(n1709), .B(n1362), .Z(n1329) );
  CENX1 U1838 ( .A(n1709), .B(b[24]), .Z(n1327) );
  CENX1 U1839 ( .A(n1712), .B(b[24]), .Z(n1294) );
  CENX1 U1840 ( .A(n1712), .B(b[25]), .Z(n1293) );
  CENX1 U1841 ( .A(n1709), .B(b[26]), .Z(n1325) );
  CENX1 U1842 ( .A(n1709), .B(b[27]), .Z(n1324) );
  CENX1 U1843 ( .A(n1708), .B(n104), .Z(n1075) );
  CENX1 U1844 ( .A(n1706), .B(n109), .Z(n1070) );
  CENX1 U1845 ( .A(n1706), .B(n104), .Z(n1077) );
  CENX1 U1846 ( .A(n1703), .B(n109), .Z(n1071) );
  CENX1 U1847 ( .A(n1710), .B(b[31]), .Z(n1320) );
  CENX1 U1848 ( .A(n1703), .B(n104), .Z(n1078) );
  CND2X1 U1849 ( .A(n100), .B(n1388), .Z(n102) );
  CEOXL U1850 ( .A(a[24]), .B(n1763), .Z(n1388) );
  CND2X2 U1851 ( .A(n1392), .B(n74), .Z(n77) );
  CNIVX1 U1852 ( .A(n116), .Z(n1703) );
  CEOXL U1853 ( .A(a[20]), .B(n1757), .Z(n1390) );
  CND2X1 U1854 ( .A(n1387), .B(n105), .Z(n107) );
  CEOXL U1855 ( .A(a[26]), .B(n104), .Z(n1387) );
  CNIVX1 U1856 ( .A(n1379), .Z(n1695) );
  CEOXL U1857 ( .A(a[22]), .B(n1761), .Z(n1389) );
  COR2X1 U1858 ( .A(n739), .B(n1568), .Z(n1561) );
  CNIVX1 U1859 ( .A(n116), .Z(n1704) );
  CND2X1 U1860 ( .A(n739), .B(n1568), .Z(n274) );
  CND2X1 U1861 ( .A(n1567), .B(n1565), .Z(n279) );
  CND2X1 U1862 ( .A(n1386), .B(n110), .Z(n112) );
  CEOXL U1863 ( .A(a[28]), .B(n109), .Z(n1386) );
  CNIVX1 U1864 ( .A(n1371), .Z(n1702) );
  CEOX1 U1865 ( .A(n1714), .B(a[4]), .Z(n1562) );
  CEOX1 U1866 ( .A(n1720), .B(a[6]), .Z(n1563) );
  CEOX1 U1867 ( .A(n1727), .B(a[8]), .Z(n1564) );
  CIVX2 U1868 ( .A(n12), .Z(n1717) );
  CND2X1 U1869 ( .A(n1385), .B(n114), .Z(n115) );
  CEOXL U1870 ( .A(a[30]), .B(a[31]), .Z(n1385) );
  CENX1 U1871 ( .A(n144), .B(n1685), .Z(n1766) );
  CND2XL U1872 ( .A(n1690), .B(n1686), .Z(n144) );
  CENX1 U1873 ( .A(n142), .B(n286), .Z(product[8]) );
  CND2XL U1874 ( .A(n1691), .B(n1689), .Z(n142) );
  CEOXL U1875 ( .A(n289), .B(n143), .Z(n1765) );
  CND2XL U1876 ( .A(n336), .B(n1687), .Z(n143) );
  CENX1 U1877 ( .A(n1715), .B(n1366), .Z(n1300) );
  CENX1 U1878 ( .A(n1721), .B(n1366), .Z(n1269) );
  CENX1 U1879 ( .A(n1728), .B(n1366), .Z(n1240) );
  CENX1 U1880 ( .A(n1735), .B(n1366), .Z(n1213) );
  CENX1 U1881 ( .A(n1740), .B(n1366), .Z(n1188) );
  CENX1 U1882 ( .A(n1725), .B(n1368), .Z(n1242) );
  CENX1 U1883 ( .A(n1716), .B(n1368), .Z(n1302) );
  CENX1 U1884 ( .A(n1736), .B(n1368), .Z(n1215) );
  CENX1 U1885 ( .A(n1744), .B(n1368), .Z(n1146) );
  CENX4 U1886 ( .A(n1710), .B(a[2]), .Z(n15) );
  CND2X4 U1887 ( .A(n1399), .B(n15), .Z(n18) );
  CND2X4 U1888 ( .A(n1395), .B(n50), .Z(n53) );
  CIVXL U1889 ( .A(n1717), .Z(n1711) );
  CIVXL U1890 ( .A(n1717), .Z(n1713) );
  CIVXL U1891 ( .A(n1717), .Z(n1714) );
  CIVXL U1892 ( .A(n1717), .Z(n1715) );
  CIVXL U1893 ( .A(n1717), .Z(n1716) );
  CIVXL U1894 ( .A(n1723), .Z(n1718) );
  CIVXL U1895 ( .A(n1723), .Z(n1719) );
  CIVXL U1896 ( .A(n1723), .Z(n1720) );
  CIVXL U1897 ( .A(n1723), .Z(n1721) );
  CIVXL U1898 ( .A(n1723), .Z(n1722) );
  CIVXL U1899 ( .A(n1730), .Z(n1724) );
  CIVXL U1900 ( .A(n1731), .Z(n1725) );
  CIVXL U1901 ( .A(n1731), .Z(n1726) );
  CIVXL U1902 ( .A(n1732), .Z(n1728) );
  CIVXL U1903 ( .A(n1732), .Z(n1729) );
  CIVXL U1904 ( .A(n30), .Z(n1730) );
  CIVXL U1905 ( .A(n30), .Z(n1731) );
  CIVXL U1906 ( .A(n30), .Z(n1732) );
  CIVXL U1907 ( .A(n1738), .Z(n1733) );
  CIVXL U1908 ( .A(n1739), .Z(n1734) );
  CIVXL U1909 ( .A(n1738), .Z(n1735) );
  CIVXL U1910 ( .A(n1739), .Z(n1736) );
  CIVXL U1911 ( .A(n1739), .Z(n1737) );
  CIVXL U1912 ( .A(n39), .Z(n1738) );
  CIVX1 U1913 ( .A(n48), .Z(n1742) );
  CIVXL U1914 ( .A(n1752), .Z(n1747) );
  CIVXL U1915 ( .A(n1752), .Z(n1748) );
  CIVXL U1916 ( .A(n1752), .Z(n1749) );
  CIVXL U1917 ( .A(n1752), .Z(n1750) );
  CIVXL U1918 ( .A(n1752), .Z(n1751) );
  CIVX1 U1919 ( .A(n71), .Z(n1752) );
  CIVXL U1920 ( .A(n1522), .Z(n1754) );
  CIVXL U1921 ( .A(n79), .Z(n1755) );
  CIVXL U1922 ( .A(n1759), .Z(n1756) );
  CIVXL U1923 ( .A(n1760), .Z(n1757) );
  CIVXL U1924 ( .A(n1760), .Z(n1758) );
  CIVXL U1925 ( .A(n86), .Z(n1759) );
  CIVXL U1926 ( .A(n86), .Z(n1760) );
  CIVX1 U1927 ( .A(n93), .Z(n1762) );
  CIVX1 U1928 ( .A(n99), .Z(n1764) );
  CIVX2 U1929 ( .A(n303), .Z(n340) );
  CIVX2 U1930 ( .A(n295), .Z(n338) );
  CIVX2 U1931 ( .A(n1688), .Z(n336) );
  CIVX2 U1932 ( .A(n265), .Z(n332) );
  CIVX2 U1933 ( .A(n262), .Z(n331) );
  CIVX2 U1934 ( .A(n251), .Z(n329) );
  CIVX2 U1935 ( .A(n224), .Z(n325) );
  CIVX2 U1936 ( .A(n159), .Z(n315) );
  CIVX2 U1937 ( .A(n151), .Z(n313) );
  CIVX2 U1938 ( .A(n312), .Z(n310) );
  CIVX2 U1939 ( .A(n309), .Z(n307) );
  CIVX2 U1940 ( .A(n301), .Z(n299) );
  CIVX2 U1941 ( .A(n1686), .Z(n291) );
  CIVX2 U1942 ( .A(n1689), .Z(n283) );
  CIVX2 U1943 ( .A(n281), .Z(n280) );
  CIVX2 U1944 ( .A(n279), .Z(n277) );
  CIVX2 U1945 ( .A(n274), .Z(n272) );
  CIVX2 U1946 ( .A(n268), .Z(n267) );
  CIVX2 U1947 ( .A(n259), .Z(n258) );
  CIVX2 U1948 ( .A(n257), .Z(n255) );
  CIVX2 U1949 ( .A(n256), .Z(n330) );
  CIVX2 U1950 ( .A(n247), .Z(n245) );
  CIVX2 U1951 ( .A(n1539), .Z(n240) );
  CIVX2 U1952 ( .A(n234), .Z(n327) );
  CIVX2 U1953 ( .A(n232), .Z(n230) );
  CIVX2 U1954 ( .A(n214), .Z(n212) );
  CIVX2 U1955 ( .A(n202), .Z(n204) );
  CIVX2 U1956 ( .A(n201), .Z(n322) );
  CIVX2 U1957 ( .A(n192), .Z(n190) );
  CIVX2 U1958 ( .A(n187), .Z(n185) );
  CIVX2 U1959 ( .A(n177), .Z(n175) );
  CIVX2 U1960 ( .A(n172), .Z(n170) );
  CIVX2 U1961 ( .A(n165), .Z(n163) );
  CIVX2 U1962 ( .A(n157), .Z(n155) );
  CIVX2 U1963 ( .A(n104), .Z(n1412) );
  CIVX2 U1964 ( .A(n109), .Z(n1411) );
endmodule


module calc_DW02_mult_2_stage_5 ( A, B, TC, CLK, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC, CLK;
  wire   n23, n24, n25, n26, n27, n28, \A_extended[32] , \B_extended[32] , n6,
         n8, n10, n12, n14, n16, n17, n18, n19, n20, n21, n22;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33;
  assign \A_extended[32]  = A[31];
  assign \B_extended[32]  = B[31];

  calc_DW_mult_tc_16 mult_96 ( .a({\A_extended[32] , \A_extended[32] , A[30:0]}), .b({\B_extended[32] , \B_extended[32] , B[30:0]}), .product({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, PRODUCT[31:6], n23, 
        n24, n25, n26, n27, n28}), .dw6_CLK(CLK) );
  CFD1QXL clk_r_REG132_S1 ( .D(n28), .CP(CLK), .Q(n17) );
  CFD1QXL clk_r_REG131_S1 ( .D(n27), .CP(CLK), .Q(n18) );
  CFD1QXL clk_r_REG125_S1 ( .D(n23), .CP(CLK), .Q(n22) );
  CFD1QXL clk_r_REG129_S1 ( .D(n25), .CP(CLK), .Q(n20) );
  CFD1QXL clk_r_REG130_S1 ( .D(n26), .CP(CLK), .Q(n19) );
  CFD1QXL clk_r_REG128_S1 ( .D(n24), .CP(CLK), .Q(n21) );
  CIVDXL U1 ( .A(n21), .Z1(n6) );
  CNIVX1 U2 ( .A(n6), .Z(PRODUCT[4]) );
  CIVDXL U3 ( .A(n19), .Z1(n8) );
  CNIVX1 U4 ( .A(n8), .Z(PRODUCT[2]) );
  CIVDXL U5 ( .A(n18), .Z1(n10) );
  CNIVX1 U6 ( .A(n10), .Z(PRODUCT[1]) );
  CIVDXL U7 ( .A(n17), .Z1(n12) );
  CNIVX1 U8 ( .A(n12), .Z(PRODUCT[0]) );
  CIVDXL U9 ( .A(n22), .Z1(n14) );
  CNIVX1 U10 ( .A(n14), .Z(PRODUCT[5]) );
  CIVDXL U11 ( .A(n20), .Z1(n16) );
  CNIVX1 U12 ( .A(n16), .Z(PRODUCT[3]) );
endmodule


module calc_DW_mult_tc_17 ( a, b, product, dw4_CLK );
  input [32:0] a;
  input [32:0] b;
  output [65:0] product;
  input dw4_CLK;
  wire   n3, n6, n9, n12, n15, n18, n21, n24, n27, n30, n33, n36, n39, n42,
         n44, n48, n50, n53, n55, n58, n61, n63, n66, n69, n71, n74, n77, n79,
         n82, n84, n86, n89, n91, n93, n95, n97, n99, n100, n102, n104, n105,
         n107, n109, n110, n112, n113, n114, n115, n116, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n155, n157,
         n158, n159, n160, n161, n163, n165, n166, n167, n168, n170, n172,
         n173, n175, n177, n178, n179, n180, n181, n182, n183, n185, n187,
         n188, n190, n192, n193, n194, n195, n197, n199, n200, n201, n202,
         n204, n207, n208, n209, n210, n212, n214, n215, n217, n219, n221,
         n222, n223, n224, n225, n226, n227, n228, n230, n232, n233, n234,
         n235, n237, n240, n241, n242, n243, n245, n247, n248, n249, n250,
         n251, n252, n253, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n272, n274, n275,
         n277, n278, n279, n280, n281, n283, n285, n286, n287, n288, n289,
         n291, n293, n294, n295, n296, n297, n299, n301, n302, n303, n304,
         n305, n307, n309, n310, n311, n312, n313, n315, n322, n325, n327,
         n329, n330, n331, n332, n334, n336, n338, n340, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1394,
         n1395, n1396, n1397, n1398, n1399, n1410, n1411, n1412, n1742, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741;
  assign n3 = a[1];
  assign n12 = a[3];
  assign n21 = a[5];
  assign n30 = a[7];
  assign n39 = a[9];
  assign n48 = a[11];
  assign n55 = a[13];
  assign n63 = a[15];
  assign n71 = a[17];
  assign n79 = a[19];
  assign n86 = a[21];
  assign n93 = a[23];
  assign n99 = a[25];
  assign n104 = a[27];
  assign n109 = a[29];
  assign n113 = a[32];
  assign n116 = b[0];
  assign n1361 = b[23];
  assign n1362 = b[22];
  assign n1363 = b[21];
  assign n1364 = b[20];
  assign n1365 = b[19];
  assign n1366 = b[18];
  assign n1367 = b[17];
  assign n1368 = b[16];
  assign n1369 = b[15];
  assign n1370 = b[14];
  assign n1371 = b[13];
  assign n1372 = b[12];
  assign n1373 = b[11];
  assign n1374 = b[10];
  assign n1375 = b[9];
  assign n1376 = b[8];
  assign n1377 = b[7];
  assign n1378 = b[6];
  assign n1379 = b[5];
  assign n1380 = b[4];
  assign n1381 = b[3];
  assign n1382 = b[2];
  assign n1383 = b[1];
  assign n1679 = dw4_CLK;

  CEO3X2 U350 ( .A(n362), .B(n344), .C(n360), .Z(n343) );
  CEO3X2 U351 ( .A(n364), .B(n346), .C(n345), .Z(n344) );
  CEO3X2 U352 ( .A(n1670), .B(n366), .C(n1671), .Z(n345) );
  CEO3X2 U353 ( .A(n1668), .B(n1669), .C(n1667), .Z(n346) );
  CEO3X2 U354 ( .A(n351), .B(n372), .C(n370), .Z(n347) );
  CEO3X2 U355 ( .A(n353), .B(n352), .C(n374), .Z(n348) );
  CEO3X2 U356 ( .A(n356), .B(n355), .C(n354), .Z(n349) );
  CEO3X2 U357 ( .A(n380), .B(n378), .C(n376), .Z(n350) );
  CEO3X2 U358 ( .A(n384), .B(n357), .C(n382), .Z(n351) );
  CEO3X2 U359 ( .A(n926), .B(n950), .C(n1034), .Z(n352) );
  CEO3X2 U360 ( .A(n850), .B(n866), .C(n1004), .Z(n353) );
  CEO3X2 U361 ( .A(n794), .B(n904), .C(n976), .Z(n354) );
  CEO3X2 U362 ( .A(n824), .B(n836), .C(n884), .Z(n355) );
  CEO3X2 U363 ( .A(n800), .B(n778), .C(n814), .Z(n356) );
  CFA1X1 U365 ( .A(n363), .B(n361), .CI(n388), .CO(n358), .S(n359) );
  CFA1X1 U366 ( .A(n367), .B(n390), .CI(n365), .CO(n360), .S(n361) );
  CFA1X1 U367 ( .A(n1666), .B(n392), .CI(n394), .CO(n362), .S(n363) );
  CFA1X1 U368 ( .A(n1662), .B(n1665), .CI(n1664), .CO(n364), .S(n365) );
  CFA1X1 U369 ( .A(n1658), .B(n1663), .CI(n1660), .CO(n366), .S(n367) );
  CFA1X1 U370 ( .A(n381), .B(n377), .CI(n379), .CO(n368), .S(n369) );
  CFA1X1 U371 ( .A(n404), .B(n402), .CI(n383), .CO(n370), .S(n371) );
  CFA1X1 U372 ( .A(n408), .B(n385), .CI(n406), .CO(n372), .S(n373) );
  CFA1X1 U373 ( .A(n927), .B(n410), .CI(n412), .CO(n374), .S(n375) );
  CFA1X1 U374 ( .A(n885), .B(n1035), .CI(n951), .CO(n376), .S(n377) );
  CFA1X1 U375 ( .A(n851), .B(n1005), .CI(n905), .CO(n378), .S(n379) );
  CFA1X1 U376 ( .A(n837), .B(n977), .CI(n867), .CO(n380), .S(n381) );
  CFA1X1 U377 ( .A(n797), .B(n825), .CI(n815), .CO(n382), .S(n383) );
  CFA1X1 U378 ( .A(n795), .B(n801), .CI(n807), .CO(n384), .S(n385) );
  CFA1X1 U379 ( .A(n391), .B(n389), .CI(n416), .CO(n386), .S(n387) );
  CFA1X1 U380 ( .A(n395), .B(n418), .CI(n393), .CO(n388), .S(n389) );
  CFA1X1 U381 ( .A(n1661), .B(n420), .CI(n422), .CO(n390), .S(n391) );
  CFA1X1 U382 ( .A(n1657), .B(n1659), .CI(n1655), .CO(n392), .S(n393) );
  CFA1X1 U383 ( .A(n1656), .B(n1653), .CI(n1651), .CO(n394), .S(n395) );
  CFA1X1 U384 ( .A(n409), .B(n405), .CI(n407), .CO(n396), .S(n397) );
  CFA1X1 U385 ( .A(n430), .B(n411), .CI(n432), .CO(n398), .S(n399) );
  CFA1X1 U386 ( .A(n438), .B(n434), .CI(n436), .CO(n400), .S(n401) );
  CFA1X1 U387 ( .A(n928), .B(n413), .CI(n952), .CO(n402), .S(n403) );
  CFA1X1 U388 ( .A(n852), .B(n1036), .CI(n886), .CO(n404), .S(n405) );
  CFA1X1 U389 ( .A(n798), .B(n1006), .CI(n906), .CO(n406), .S(n407) );
  CFA1X1 U390 ( .A(n838), .B(n978), .CI(n868), .CO(n408), .S(n409) );
  CFA1X1 U391 ( .A(n802), .B(n826), .CI(n816), .CO(n410), .S(n411) );
  CHA1X1 U392 ( .A(n808), .B(n779), .CO(n412), .S(n413) );
  CFA1X1 U393 ( .A(n419), .B(n417), .CI(n442), .CO(n414), .S(n415) );
  CFA1X1 U394 ( .A(n423), .B(n444), .CI(n421), .CO(n416), .S(n417) );
  CFA1X1 U395 ( .A(n1654), .B(n446), .CI(n1648), .CO(n418), .S(n419) );
  CFA1X1 U396 ( .A(n1646), .B(n1652), .CI(n1650), .CO(n420), .S(n421) );
  CFA1X1 U397 ( .A(n1649), .B(n1644), .CI(n1642), .CO(n422), .S(n423) );
  CFA1X1 U398 ( .A(n437), .B(n433), .CI(n435), .CO(n424), .S(n425) );
  CFA1X1 U399 ( .A(n460), .B(n456), .CI(n439), .CO(n426), .S(n427) );
  CFA1X1 U400 ( .A(n464), .B(n458), .CI(n462), .CO(n428), .S(n429) );
  CFA1X1 U401 ( .A(n887), .B(n953), .CI(n929), .CO(n430), .S(n431) );
  CFA1X1 U402 ( .A(n869), .B(n1007), .CI(n1037), .CO(n432), .S(n433) );
  CFA1X1 U403 ( .A(n853), .B(n979), .CI(n907), .CO(n434), .S(n435) );
  CFA1X1 U404 ( .A(n817), .B(n839), .CI(n827), .CO(n436), .S(n437) );
  CFA1X1 U405 ( .A(n799), .B(n803), .CI(n809), .CO(n438), .S(n439) );
  CFA1X1 U406 ( .A(n445), .B(n443), .CI(n468), .CO(n440), .S(n441) );
  CFA1X1 U407 ( .A(n1647), .B(n470), .CI(n447), .CO(n442), .S(n443) );
  CFA1X1 U408 ( .A(n1640), .B(n472), .CI(n1645), .CO(n444), .S(n445) );
  CFA1X1 U409 ( .A(n1641), .B(n1643), .CI(n1638), .CO(n446), .S(n447) );
  CFA1X1 U410 ( .A(n459), .B(n478), .CI(n457), .CO(n448), .S(n449) );
  CFA1X1 U411 ( .A(n480), .B(n461), .CI(n463), .CO(n450), .S(n451) );
  CFA1X1 U412 ( .A(n486), .B(n482), .CI(n484), .CO(n452), .S(n453) );
  CFA1X1 U413 ( .A(n930), .B(n488), .CI(n465), .CO(n454), .S(n455) );
  CFA1X1 U414 ( .A(n870), .B(n1038), .CI(n954), .CO(n456), .S(n457) );
  CFA1X1 U415 ( .A(n854), .B(n980), .CI(n888), .CO(n458), .S(n459) );
  CFA1X1 U416 ( .A(n804), .B(n1008), .CI(n908), .CO(n460), .S(n461) );
  CFA1X1 U417 ( .A(n780), .B(n840), .CI(n828), .CO(n462), .S(n463) );
  CHA1X1 U418 ( .A(n810), .B(n818), .CO(n464), .S(n465) );
  CFA1X1 U419 ( .A(n471), .B(n469), .CI(n492), .CO(n466), .S(n467) );
  CFA1X1 U420 ( .A(n496), .B(n494), .CI(n473), .CO(n468), .S(n469) );
  CFA1X1 U421 ( .A(n1635), .B(n1639), .CI(n1637), .CO(n470), .S(n471) );
  CFA1X1 U422 ( .A(n1631), .B(n1636), .CI(n1633), .CO(n472), .S(n473) );
  CFA1X1 U423 ( .A(n485), .B(n481), .CI(n483), .CO(n474), .S(n475) );
  CFA1X1 U424 ( .A(n508), .B(n487), .CI(n504), .CO(n476), .S(n477) );
  CFA1X1 U425 ( .A(n510), .B(n489), .CI(n506), .CO(n478), .S(n479) );
  CFA1X1 U426 ( .A(n931), .B(n512), .CI(n955), .CO(n480), .S(n481) );
  CFA1X1 U427 ( .A(n871), .B(n981), .CI(n1039), .CO(n482), .S(n483) );
  CFA1X1 U428 ( .A(n855), .B(n1009), .CI(n909), .CO(n484), .S(n485) );
  CFA1X1 U429 ( .A(n829), .B(n889), .CI(n841), .CO(n486), .S(n487) );
  CFA1X1 U430 ( .A(n805), .B(n819), .CI(n811), .CO(n488), .S(n489) );
  CFA1X1 U431 ( .A(n495), .B(n493), .CI(n516), .CO(n490), .S(n491) );
  CFA1X1 U432 ( .A(n520), .B(n518), .CI(n497), .CO(n492), .S(n493) );
  CFA1X1 U433 ( .A(n1629), .B(n1634), .CI(n1632), .CO(n494), .S(n495) );
  CFA1X1 U434 ( .A(n1625), .B(n1630), .CI(n1627), .CO(n496), .S(n497) );
  CFA1X1 U435 ( .A(n509), .B(n505), .CI(n507), .CO(n498), .S(n499) );
  CFA1X1 U436 ( .A(n530), .B(n511), .CI(n528), .CO(n500), .S(n501) );
  CFA1X1 U437 ( .A(n513), .B(n532), .CI(n534), .CO(n502), .S(n503) );
  CFA1X1 U438 ( .A(n932), .B(n1040), .CI(n956), .CO(n504), .S(n505) );
  CFA1X1 U439 ( .A(n856), .B(n982), .CI(n872), .CO(n506), .S(n507) );
  CFA1X1 U440 ( .A(n812), .B(n1010), .CI(n910), .CO(n508), .S(n509) );
  CFA1X1 U441 ( .A(n830), .B(n890), .CI(n842), .CO(n510), .S(n511) );
  CHA1X1 U442 ( .A(n781), .B(n820), .CO(n512), .S(n513) );
  CFA1X1 U443 ( .A(n519), .B(n517), .CI(n538), .CO(n514), .S(n515) );
  CFA1X1 U444 ( .A(n542), .B(n521), .CI(n540), .CO(n516), .S(n517) );
  CFA1X1 U445 ( .A(n1622), .B(n1628), .CI(n1626), .CO(n518), .S(n519) );
  CFA1X1 U446 ( .A(n1623), .B(n1624), .CI(n1620), .CO(n520), .S(n521) );
  CFA1X1 U447 ( .A(n533), .B(n548), .CI(n531), .CO(n522), .S(n523) );
  CFA1X1 U448 ( .A(n550), .B(n535), .CI(n552), .CO(n524), .S(n525) );
  CFA1X1 U449 ( .A(n933), .B(n554), .CI(n556), .CO(n526), .S(n527) );
  CFA1X1 U450 ( .A(n891), .B(n1041), .CI(n957), .CO(n528), .S(n529) );
  CFA1X1 U451 ( .A(n857), .B(n1011), .CI(n911), .CO(n530), .S(n531) );
  CFA1X1 U452 ( .A(n843), .B(n983), .CI(n873), .CO(n532), .S(n533) );
  CFA1X1 U453 ( .A(n813), .B(n831), .CI(n821), .CO(n534), .S(n535) );
  CFA1X1 U454 ( .A(n541), .B(n539), .CI(n560), .CO(n536), .S(n537) );
  CFA1X1 U455 ( .A(n1621), .B(n562), .CI(n543), .CO(n538), .S(n539) );
  CFA1X1 U456 ( .A(n1614), .B(n1616), .CI(n1619), .CO(n540), .S(n541) );
  CFA1X1 U457 ( .A(n1617), .B(n1612), .CI(n1618), .CO(n542), .S(n543) );
  CFA1X1 U458 ( .A(n572), .B(n553), .CI(n555), .CO(n544), .S(n545) );
  CFA1X1 U459 ( .A(n576), .B(n570), .CI(n574), .CO(n546), .S(n547) );
  CFA1X1 U460 ( .A(n934), .B(n557), .CI(n958), .CO(n548), .S(n549) );
  CFA1X1 U461 ( .A(n858), .B(n1042), .CI(n892), .CO(n550), .S(n551) );
  CFA1X1 U462 ( .A(n822), .B(n984), .CI(n912), .CO(n552), .S(n553) );
  CFA1X1 U463 ( .A(n844), .B(n1012), .CI(n874), .CO(n554), .S(n555) );
  CHA1X1 U464 ( .A(n782), .B(n832), .CO(n556), .S(n557) );
  CFA1X1 U465 ( .A(n563), .B(n561), .CI(n580), .CO(n558), .S(n559) );
  CFA1X1 U466 ( .A(n1613), .B(n582), .CI(n1615), .CO(n560), .S(n561) );
  CFA1X1 U467 ( .A(n1608), .B(n1610), .CI(n1611), .CO(n562), .S(n563) );
  CFA1X1 U468 ( .A(n573), .B(n588), .CI(n571), .CO(n564), .S(n565) );
  CFA1X1 U469 ( .A(n590), .B(n575), .CI(n577), .CO(n566), .S(n567) );
  CFA1X1 U470 ( .A(n596), .B(n594), .CI(n592), .CO(n568), .S(n569) );
  CFA1X1 U471 ( .A(n893), .B(n959), .CI(n935), .CO(n570), .S(n571) );
  CFA1X1 U472 ( .A(n875), .B(n1013), .CI(n1043), .CO(n572), .S(n573) );
  CFA1X1 U473 ( .A(n859), .B(n985), .CI(n913), .CO(n574), .S(n575) );
  CFA1X1 U475 ( .A(n583), .B(n581), .CI(n600), .CO(n578), .S(n579) );
  CFA1X1 U476 ( .A(n1607), .B(n602), .CI(n1609), .CO(n580), .S(n581) );
  CFA1X1 U477 ( .A(n1603), .B(n1605), .CI(n1606), .CO(n582), .S(n583) );
  CFA1X1 U478 ( .A(n595), .B(n591), .CI(n593), .CO(n584), .S(n585) );
  CFA1X1 U479 ( .A(n610), .B(n608), .CI(n612), .CO(n586), .S(n587) );
  CFA1X1 U480 ( .A(n936), .B(n614), .CI(n597), .CO(n588), .S(n589) );
  CFA1X1 U481 ( .A(n876), .B(n1044), .CI(n960), .CO(n590), .S(n591) );
  CFA1X1 U482 ( .A(n860), .B(n1014), .CI(n894), .CO(n592), .S(n593) );
  CFA1X1 U483 ( .A(n834), .B(n986), .CI(n914), .CO(n594), .S(n595) );
  CHA1X1 U484 ( .A(n783), .B(n846), .CO(n596), .S(n597) );
  CFA1X1 U485 ( .A(n603), .B(n601), .CI(n618), .CO(n598), .S(n599) );
  CFA1X1 U486 ( .A(n1602), .B(n1600), .CI(n1604), .CO(n600), .S(n601) );
  CFA1X1 U487 ( .A(n1601), .B(n1598), .CI(n1596), .CO(n602), .S(n603) );
  CFA1X1 U488 ( .A(n615), .B(n611), .CI(n613), .CO(n604), .S(n605) );
  CFA1X1 U489 ( .A(n630), .B(n626), .CI(n628), .CO(n606), .S(n607) );
  CFA1X1 U490 ( .A(n915), .B(n632), .CI(n937), .CO(n608), .S(n609) );
  CFA1X1 U491 ( .A(n895), .B(n1015), .CI(n961), .CO(n610), .S(n611) );
  CFA1X1 U492 ( .A(n877), .B(n987), .CI(n1045), .CO(n612), .S(n613) );
  CFA1X1 U493 ( .A(n835), .B(n861), .CI(n847), .CO(n614), .S(n615) );
  CFA1X1 U494 ( .A(n1599), .B(n619), .CI(n636), .CO(n616), .S(n617) );
  CFA1X1 U495 ( .A(n1595), .B(n638), .CI(n1597), .CO(n618), .S(n619) );
  CFA1X1 U496 ( .A(n627), .B(n640), .CI(n642), .CO(n620), .S(n621) );
  CFA1X1 U497 ( .A(n646), .B(n629), .CI(n631), .CO(n622), .S(n623) );
  CFA1X1 U498 ( .A(n633), .B(n644), .CI(n648), .CO(n624), .S(n625) );
  CFA1X1 U499 ( .A(n896), .B(n1046), .CI(n962), .CO(n626), .S(n627) );
  CFA1X1 U500 ( .A(n848), .B(n1016), .CI(n938), .CO(n628), .S(n629) );
  CFA1X1 U501 ( .A(n862), .B(n988), .CI(n916), .CO(n630), .S(n631) );
  CHA1X1 U502 ( .A(n784), .B(n878), .CO(n632), .S(n633) );
  CFA1X1 U503 ( .A(n639), .B(n637), .CI(n652), .CO(n634), .S(n635) );
  CFA1X1 U504 ( .A(n1593), .B(n1591), .CI(n1594), .CO(n636), .S(n637) );
  CFA1X1 U505 ( .A(n1592), .B(n1589), .CI(n1587), .CO(n638), .S(n639) );
  CFA1X1 U506 ( .A(n662), .B(n647), .CI(n649), .CO(n640), .S(n641) );
  CFA1X1 U507 ( .A(n939), .B(n660), .CI(n664), .CO(n642), .S(n643) );
  CFA1X1 U508 ( .A(n917), .B(n1047), .CI(n963), .CO(n644), .S(n645) );
  CFA1X1 U509 ( .A(n897), .B(n1017), .CI(n989), .CO(n646), .S(n647) );
  CFA1X1 U510 ( .A(n849), .B(n879), .CI(n863), .CO(n648), .S(n649) );
  CFA1X1 U511 ( .A(n1590), .B(n653), .CI(n668), .CO(n650), .S(n651) );
  CFA1X1 U512 ( .A(n1586), .B(n1585), .CI(n1588), .CO(n652), .S(n653) );
  CFA1X1 U513 ( .A(n663), .B(n672), .CI(n661), .CO(n654), .S(n655) );
  CFA1X1 U514 ( .A(n678), .B(n674), .CI(n676), .CO(n656), .S(n657) );
  CFA1X1 U515 ( .A(n864), .B(n665), .CI(n918), .CO(n658), .S(n659) );
  CFA1X1 U516 ( .A(n898), .B(n990), .CI(n964), .CO(n660), .S(n661) );
  CFA1X1 U517 ( .A(n880), .B(n1018), .CI(n1048), .CO(n662), .S(n663) );
  CHA1X1 U518 ( .A(n785), .B(n940), .CO(n664), .S(n665) );
  CFA1X1 U519 ( .A(n1584), .B(n669), .CI(n682), .CO(n666), .S(n667) );
  CFA1X1 U520 ( .A(n1580), .B(n1582), .CI(n1583), .CO(n668), .S(n669) );
  CFA1X1 U521 ( .A(n679), .B(n675), .CI(n677), .CO(n670), .S(n671) );
  CFA1X1 U522 ( .A(n692), .B(n690), .CI(n688), .CO(n672), .S(n673) );
  CFA1X1 U523 ( .A(n941), .B(n1049), .CI(n965), .CO(n674), .S(n675) );
  CFA1X1 U524 ( .A(n919), .B(n1019), .CI(n991), .CO(n676), .S(n677) );
  CFA1X1 U525 ( .A(n865), .B(n899), .CI(n881), .CO(n678), .S(n679) );
  CFA1X1 U526 ( .A(n1581), .B(n683), .CI(n696), .CO(n680), .S(n681) );
  CFA1X1 U527 ( .A(n1576), .B(n1579), .CI(n1578), .CO(n682), .S(n683) );
  CFA1X1 U528 ( .A(n702), .B(n689), .CI(n691), .CO(n684), .S(n685) );
  CFA1X1 U529 ( .A(n920), .B(n704), .CI(n693), .CO(n686), .S(n687) );
  CFA1X1 U530 ( .A(n882), .B(n966), .CI(n942), .CO(n688), .S(n689) );
  CFA1X1 U531 ( .A(n900), .B(n992), .CI(n1050), .CO(n690), .S(n691) );
  CHA1X1 U532 ( .A(n786), .B(n1020), .CO(n692), .S(n693) );
  CFA1X1 U533 ( .A(n1577), .B(n697), .CI(n708), .CO(n694), .S(n695) );
  CFA1X1 U534 ( .A(n1574), .B(n1573), .CI(n1575), .CO(n696), .S(n697) );
  CFA1X1 U535 ( .A(n712), .B(n705), .CI(n714), .CO(n698), .S(n699) );
  CFA1X1 U536 ( .A(n967), .B(n716), .CI(n1051), .CO(n700), .S(n701) );
  CFA1X1 U537 ( .A(n943), .B(n993), .CI(n1021), .CO(n702), .S(n703) );
  CFA1X1 U538 ( .A(n883), .B(n921), .CI(n901), .CO(n704), .S(n705) );
  CFA1X1 U539 ( .A(n1572), .B(n709), .CI(n1569), .CO(n706), .S(n707) );
  CFA1X1 U540 ( .A(n1570), .B(n1567), .CI(n1571), .CO(n708), .S(n709) );
  CFA1X1 U541 ( .A(n717), .B(n724), .CI(n726), .CO(n710), .S(n711) );
  CFA1X1 U542 ( .A(n922), .B(n968), .CI(n944), .CO(n712), .S(n713) );
  CFA1X1 U543 ( .A(n902), .B(n994), .CI(n1052), .CO(n714), .S(n715) );
  CHA1X1 U544 ( .A(n787), .B(n1022), .CO(n716), .S(n717) );
  CFA1X1 U545 ( .A(n1565), .B(n1568), .CI(n1566), .CO(n718), .S(n719) );
  CFA1X1 U546 ( .A(n727), .B(n732), .CI(n725), .CO(n720), .S(n721) );
  CFA1X1 U547 ( .A(n1053), .B(n734), .CI(n736), .CO(n722), .S(n723) );
  CFA1X1 U548 ( .A(n969), .B(n1023), .CI(n995), .CO(n724), .S(n725) );
  CFA1X1 U549 ( .A(n903), .B(n945), .CI(n923), .CO(n726), .S(n727) );
  CFA1X1 U550 ( .A(n1563), .B(n1564), .CI(n1562), .CO(n728), .S(n729) );
  CFA1X1 U551 ( .A(n744), .B(n735), .CI(n742), .CO(n730), .S(n731) );
  CFA1X1 U552 ( .A(n946), .B(n737), .CI(n970), .CO(n732), .S(n733) );
  CFA1X1 U553 ( .A(n924), .B(n996), .CI(n1054), .CO(n734), .S(n735) );
  CHA1X1 U554 ( .A(n788), .B(n1024), .CO(n736), .S(n737) );
  CFA1X1 U555 ( .A(n1560), .B(n1561), .CI(n1558), .CO(n738), .S(n739) );
  CFA1X1 U556 ( .A(n752), .B(n745), .CI(n750), .CO(n740), .S(n741) );
  CFA1X1 U557 ( .A(n1055), .B(n1025), .CI(n997), .CO(n742), .S(n743) );
  CFA1X1 U558 ( .A(n925), .B(n971), .CI(n947), .CO(n744), .S(n745) );
  CFA1X1 U559 ( .A(n756), .B(n749), .CI(n751), .CO(n746), .S(n747) );
  CFA1X1 U560 ( .A(n972), .B(n758), .CI(n753), .CO(n748), .S(n749) );
  CFA1X1 U561 ( .A(n948), .B(n998), .CI(n1056), .CO(n750), .S(n751) );
  CFA1X1 U563 ( .A(n762), .B(n757), .CI(n759), .CO(n754), .S(n755) );
  CFA1X1 U564 ( .A(n1027), .B(n764), .CI(n999), .CO(n756), .S(n757) );
  CFA1X1 U565 ( .A(n949), .B(n1057), .CI(n973), .CO(n758), .S(n759) );
  CFA1X1 U566 ( .A(n765), .B(n763), .CI(n768), .CO(n760), .S(n761) );
  CFA1X1 U567 ( .A(n974), .B(n1000), .CI(n1058), .CO(n762), .S(n763) );
  CHA1X1 U568 ( .A(n790), .B(n1028), .CO(n764), .S(n765) );
  CFA1X1 U569 ( .A(n1001), .B(n769), .CI(n772), .CO(n766), .S(n767) );
  CFA1X1 U570 ( .A(n975), .B(n1029), .CI(n1059), .CO(n768), .S(n769) );
  CFA1X1 U571 ( .A(n1030), .B(n773), .CI(n1002), .CO(n770), .S(n771) );
  CHA1X1 U572 ( .A(n1060), .B(n791), .CO(n772), .S(n773) );
  CFA1X1 U573 ( .A(n1003), .B(n1031), .CI(n1061), .CO(n774), .S(n775) );
  CHA1X1 U574 ( .A(n1062), .B(n1032), .CO(n776), .S(n777) );
  COND2X1 U576 ( .A(n1066), .B(n115), .C(n114), .D(n1065), .Z(n794) );
  COND2X1 U581 ( .A(n1072), .B(n110), .C(n1411), .D(n112), .Z(n779) );
  COND2X1 U582 ( .A(n112), .B(n1069), .C(n110), .D(n1068), .Z(n796) );
  COND2X1 U583 ( .A(n112), .B(n1070), .C(n110), .D(n1069), .Z(n797) );
  COND2X1 U584 ( .A(n1071), .B(n112), .C(n110), .D(n1070), .Z(n798) );
  COND2X1 U591 ( .A(n1079), .B(n105), .C(n1412), .D(n107), .Z(n780) );
  COND2X1 U592 ( .A(n107), .B(n1074), .C(n105), .D(n1073), .Z(n800) );
  COND2X1 U593 ( .A(n1075), .B(n107), .C(n105), .D(n1074), .Z(n801) );
  COND2X1 U594 ( .A(n1076), .B(n107), .C(n105), .D(n1075), .Z(n802) );
  COND2X1 U596 ( .A(n1078), .B(n107), .C(n105), .D(n1077), .Z(n804) );
  CND2IX1 U604 ( .B(n1685), .A(n104), .Z(n1079) );
  COND2X1 U605 ( .A(n1088), .B(n100), .C(n1741), .D(n102), .Z(n781) );
  COND2X1 U607 ( .A(n102), .B(n1082), .C(n100), .D(n1081), .Z(n807) );
  COND2X1 U608 ( .A(n102), .B(n1083), .C(n100), .D(n1082), .Z(n808) );
  COND2X1 U609 ( .A(n102), .B(n1084), .C(n100), .D(n1083), .Z(n809) );
  COND2X1 U610 ( .A(n102), .B(n1085), .C(n100), .D(n1084), .Z(n810) );
  COND2X1 U611 ( .A(n102), .B(n1086), .C(n100), .D(n1085), .Z(n811) );
  COND2X1 U612 ( .A(n1087), .B(n102), .C(n100), .D(n1086), .Z(n812) );
  CND2IX1 U622 ( .B(n1685), .A(n1740), .Z(n1088) );
  COND2X1 U623 ( .A(n97), .B(n1739), .C(n95), .D(n1099), .Z(n782) );
  COND2X1 U624 ( .A(n97), .B(n1090), .C(n1089), .D(n95), .Z(n814) );
  COND2X1 U625 ( .A(n97), .B(n1091), .C(n1090), .D(n95), .Z(n815) );
  COND2X1 U626 ( .A(n97), .B(n1092), .C(n1091), .D(n95), .Z(n816) );
  COND2X1 U627 ( .A(n97), .B(n1093), .C(n1092), .D(n95), .Z(n817) );
  COND2X1 U628 ( .A(n97), .B(n1094), .C(n95), .D(n1093), .Z(n818) );
  COND2X1 U629 ( .A(n97), .B(n1095), .C(n95), .D(n1094), .Z(n819) );
  COND2X1 U630 ( .A(n97), .B(n1096), .C(n95), .D(n1095), .Z(n820) );
  COND2X1 U631 ( .A(n97), .B(n1097), .C(n95), .D(n1096), .Z(n821) );
  COND2X1 U632 ( .A(n1098), .B(n97), .C(n95), .D(n1097), .Z(n822) );
  CND2IX1 U644 ( .B(n1685), .A(n1738), .Z(n1099) );
  CND2IX1 U670 ( .B(n1685), .A(n1733), .Z(n1112) );
  COND2X1 U671 ( .A(n84), .B(n1522), .C(n82), .D(n1127), .Z(n784) );
  COND2X1 U672 ( .A(n84), .B(n1114), .C(n1113), .D(n82), .Z(n836) );
  COND2X1 U673 ( .A(n84), .B(n1115), .C(n1114), .D(n82), .Z(n837) );
  COND2X1 U674 ( .A(n84), .B(n1116), .C(n1115), .D(n82), .Z(n838) );
  COND2X1 U675 ( .A(n84), .B(n1117), .C(n1116), .D(n82), .Z(n839) );
  COND2X1 U676 ( .A(n84), .B(n1118), .C(n1117), .D(n82), .Z(n840) );
  COND2X1 U677 ( .A(n84), .B(n1119), .C(n1118), .D(n82), .Z(n841) );
  COND2X1 U678 ( .A(n84), .B(n1120), .C(n1119), .D(n82), .Z(n842) );
  COND2X1 U679 ( .A(n84), .B(n1121), .C(n1120), .D(n82), .Z(n843) );
  COND2X1 U680 ( .A(n84), .B(n1122), .C(n1121), .D(n82), .Z(n844) );
  COND2X1 U681 ( .A(n84), .B(n1123), .C(n1122), .D(n82), .Z(n845) );
  COND2X1 U682 ( .A(n84), .B(n1124), .C(n1123), .D(n82), .Z(n846) );
  COND2X1 U684 ( .A(n1126), .B(n84), .C(n1125), .D(n82), .Z(n848) );
  CND2IX1 U700 ( .B(n1685), .A(n1523), .Z(n1127) );
  COND2X1 U701 ( .A(n77), .B(n1528), .C(n74), .D(n1144), .Z(n785) );
  COND2X1 U702 ( .A(n77), .B(n1129), .C(n1128), .D(n74), .Z(n850) );
  COND2X1 U703 ( .A(n77), .B(n1130), .C(n1129), .D(n74), .Z(n851) );
  COND2X1 U704 ( .A(n77), .B(n1131), .C(n1130), .D(n74), .Z(n852) );
  COND2X1 U705 ( .A(n77), .B(n1132), .C(n1131), .D(n74), .Z(n853) );
  COND2X1 U706 ( .A(n77), .B(n1133), .C(n1132), .D(n74), .Z(n854) );
  COND2X1 U707 ( .A(n77), .B(n1134), .C(n1133), .D(n74), .Z(n855) );
  COND2X1 U708 ( .A(n77), .B(n1135), .C(n1134), .D(n74), .Z(n856) );
  COND2X1 U709 ( .A(n77), .B(n1136), .C(n1135), .D(n74), .Z(n857) );
  COND2X1 U710 ( .A(n77), .B(n1137), .C(n1136), .D(n74), .Z(n858) );
  COND2X1 U711 ( .A(n77), .B(n1138), .C(n1137), .D(n74), .Z(n859) );
  COND2X1 U712 ( .A(n77), .B(n1139), .C(n1138), .D(n74), .Z(n860) );
  COND2X1 U713 ( .A(n77), .B(n1140), .C(n1139), .D(n74), .Z(n861) );
  COND2X1 U714 ( .A(n77), .B(n1141), .C(n1140), .D(n74), .Z(n862) );
  COND2X1 U715 ( .A(n77), .B(n1142), .C(n1141), .D(n74), .Z(n863) );
  COND2X1 U716 ( .A(n77), .B(n1143), .C(n1142), .D(n74), .Z(n864) );
  CND2IX1 U734 ( .B(n1685), .A(n1728), .Z(n1144) );
  COND2X1 U737 ( .A(n69), .B(n1147), .C(n1146), .D(n66), .Z(n867) );
  COND2X1 U738 ( .A(n69), .B(n1148), .C(n1147), .D(n66), .Z(n868) );
  COND2X1 U742 ( .A(n69), .B(n1152), .C(n1151), .D(n66), .Z(n872) );
  COND2X1 U743 ( .A(n69), .B(n1153), .C(n1152), .D(n66), .Z(n873) );
  COND2X1 U745 ( .A(n69), .B(n1155), .C(n1154), .D(n66), .Z(n875) );
  COND2X1 U749 ( .A(n69), .B(n1159), .C(n1158), .D(n66), .Z(n879) );
  COND2X1 U750 ( .A(n69), .B(n1160), .C(n1159), .D(n66), .Z(n880) );
  COND2X1 U752 ( .A(n69), .B(n1162), .C(n1161), .D(n66), .Z(n882) );
  COND2X1 U773 ( .A(n61), .B(n1724), .C(n1184), .D(n58), .Z(n787) );
  COND2X1 U774 ( .A(n61), .B(n1165), .C(n1164), .D(n58), .Z(n884) );
  COND2X1 U775 ( .A(n61), .B(n1166), .C(n1165), .D(n58), .Z(n885) );
  COND2X1 U776 ( .A(n61), .B(n1167), .C(n1166), .D(n58), .Z(n886) );
  COND2X1 U777 ( .A(n61), .B(n1168), .C(n1167), .D(n58), .Z(n887) );
  COND2X1 U778 ( .A(n61), .B(n1169), .C(n1168), .D(n58), .Z(n888) );
  COND2X1 U779 ( .A(n61), .B(n1170), .C(n1169), .D(n58), .Z(n889) );
  COND2X1 U780 ( .A(n61), .B(n1171), .C(n1170), .D(n58), .Z(n890) );
  COND2X1 U781 ( .A(n61), .B(n1172), .C(n1171), .D(n58), .Z(n891) );
  COND2X1 U782 ( .A(n61), .B(n1173), .C(n1172), .D(n58), .Z(n892) );
  COND2X1 U783 ( .A(n61), .B(n1174), .C(n1173), .D(n58), .Z(n893) );
  COND2X1 U784 ( .A(n61), .B(n1175), .C(n1174), .D(n58), .Z(n894) );
  COND2X1 U785 ( .A(n61), .B(n1176), .C(n1175), .D(n58), .Z(n895) );
  COND2X1 U786 ( .A(n61), .B(n1177), .C(n1176), .D(n58), .Z(n896) );
  COND2X1 U787 ( .A(n61), .B(n1178), .C(n1177), .D(n58), .Z(n897) );
  COND2X1 U788 ( .A(n61), .B(n1179), .C(n1178), .D(n58), .Z(n898) );
  COND2X1 U789 ( .A(n61), .B(n1180), .C(n1179), .D(n58), .Z(n899) );
  COND2X1 U790 ( .A(n61), .B(n1181), .C(n1180), .D(n58), .Z(n900) );
  COND2X1 U791 ( .A(n61), .B(n1182), .C(n1181), .D(n58), .Z(n901) );
  COND2X1 U792 ( .A(n61), .B(n1183), .C(n1182), .D(n58), .Z(n902) );
  CND2IX1 U814 ( .B(n1685), .A(n1723), .Z(n1184) );
  COND2X1 U815 ( .A(n53), .B(n1721), .C(n1207), .D(n50), .Z(n788) );
  COND2X1 U816 ( .A(n53), .B(n1186), .C(n1185), .D(n50), .Z(n904) );
  COND2X1 U817 ( .A(n53), .B(n1187), .C(n1186), .D(n50), .Z(n905) );
  COND2X1 U818 ( .A(n53), .B(n1188), .C(n1187), .D(n50), .Z(n906) );
  COND2X1 U819 ( .A(n53), .B(n1189), .C(n1188), .D(n50), .Z(n907) );
  COND2X1 U820 ( .A(n53), .B(n1190), .C(n1189), .D(n50), .Z(n908) );
  COND2X1 U821 ( .A(n53), .B(n1191), .C(n1190), .D(n50), .Z(n909) );
  COND2X1 U822 ( .A(n53), .B(n1192), .C(n1191), .D(n50), .Z(n910) );
  COND2X1 U823 ( .A(n53), .B(n1193), .C(n1192), .D(n50), .Z(n911) );
  COND2X1 U824 ( .A(n53), .B(n1194), .C(n1193), .D(n50), .Z(n912) );
  COND2X1 U825 ( .A(n53), .B(n1195), .C(n1194), .D(n50), .Z(n913) );
  COND2X1 U826 ( .A(n53), .B(n1196), .C(n1195), .D(n50), .Z(n914) );
  COND2X1 U827 ( .A(n53), .B(n1197), .C(n1196), .D(n50), .Z(n915) );
  COND2X1 U828 ( .A(n53), .B(n1198), .C(n1197), .D(n50), .Z(n916) );
  COND2X1 U829 ( .A(n53), .B(n1199), .C(n1198), .D(n50), .Z(n917) );
  COND2X1 U831 ( .A(n53), .B(n1201), .C(n1200), .D(n50), .Z(n919) );
  COND2X1 U832 ( .A(n53), .B(n1202), .C(n1201), .D(n50), .Z(n920) );
  COND2X1 U834 ( .A(n53), .B(n1204), .C(n1203), .D(n50), .Z(n922) );
  COND2X1 U835 ( .A(n53), .B(n1205), .C(n1204), .D(n50), .Z(n923) );
  COND2X1 U836 ( .A(n53), .B(n1206), .C(n1205), .D(n50), .Z(n924) );
  CND2IX1 U860 ( .B(n1685), .A(n1720), .Z(n1207) );
  COND2X1 U862 ( .A(n44), .B(n1209), .C(n1208), .D(n42), .Z(n926) );
  COND2X1 U863 ( .A(n44), .B(n1210), .C(n1209), .D(n42), .Z(n927) );
  COND2X1 U864 ( .A(n44), .B(n1211), .C(n1210), .D(n42), .Z(n928) );
  COND2X1 U865 ( .A(n44), .B(n1212), .C(n1211), .D(n42), .Z(n929) );
  COND2X1 U866 ( .A(n44), .B(n1213), .C(n1212), .D(n42), .Z(n930) );
  COND2X1 U867 ( .A(n44), .B(n1214), .C(n1213), .D(n42), .Z(n931) );
  COND2X1 U868 ( .A(n44), .B(n1215), .C(n1214), .D(n42), .Z(n932) );
  COND2X1 U869 ( .A(n44), .B(n1216), .C(n1215), .D(n42), .Z(n933) );
  COND2X1 U870 ( .A(n44), .B(n1217), .C(n1216), .D(n42), .Z(n934) );
  COND2X1 U871 ( .A(n44), .B(n1218), .C(n1217), .D(n42), .Z(n935) );
  COND2X1 U872 ( .A(n44), .B(n1219), .C(n1218), .D(n42), .Z(n936) );
  COND2X1 U873 ( .A(n44), .B(n1220), .C(n1219), .D(n42), .Z(n937) );
  COND2X1 U874 ( .A(n44), .B(n1221), .C(n1220), .D(n42), .Z(n938) );
  COND2X1 U875 ( .A(n44), .B(n1222), .C(n1221), .D(n42), .Z(n939) );
  COND2X1 U877 ( .A(n44), .B(n1224), .C(n1223), .D(n42), .Z(n941) );
  COND2X1 U878 ( .A(n44), .B(n1225), .C(n1224), .D(n42), .Z(n942) );
  COND2X1 U879 ( .A(n44), .B(n1226), .C(n1225), .D(n42), .Z(n943) );
  COND2X1 U880 ( .A(n44), .B(n1227), .C(n1226), .D(n42), .Z(n944) );
  COND2X1 U881 ( .A(n44), .B(n1228), .C(n1227), .D(n42), .Z(n945) );
  COND2X1 U882 ( .A(n44), .B(n1229), .C(n1228), .D(n42), .Z(n946) );
  COND2X1 U884 ( .A(n44), .B(n1231), .C(n1230), .D(n42), .Z(n948) );
  CND2IX1 U910 ( .B(n1685), .A(n1711), .Z(n1232) );
  COND2X1 U911 ( .A(n36), .B(n1708), .C(n1259), .D(n33), .Z(n790) );
  COND2X1 U912 ( .A(n36), .B(n1234), .C(n1233), .D(n33), .Z(n950) );
  COND2X1 U913 ( .A(n36), .B(n1235), .C(n1234), .D(n33), .Z(n951) );
  COND2X1 U914 ( .A(n36), .B(n1236), .C(n1235), .D(n33), .Z(n952) );
  COND2X1 U915 ( .A(n36), .B(n1237), .C(n1236), .D(n33), .Z(n953) );
  COND2X1 U916 ( .A(n36), .B(n1238), .C(n1237), .D(n33), .Z(n954) );
  COND2X1 U917 ( .A(n36), .B(n1239), .C(n1238), .D(n33), .Z(n955) );
  COND2X1 U918 ( .A(n36), .B(n1240), .C(n1239), .D(n33), .Z(n956) );
  COND2X1 U919 ( .A(n36), .B(n1241), .C(n1240), .D(n33), .Z(n957) );
  COND2X1 U920 ( .A(n36), .B(n1242), .C(n1241), .D(n33), .Z(n958) );
  COND2X1 U921 ( .A(n36), .B(n1243), .C(n1242), .D(n33), .Z(n959) );
  COND2X1 U922 ( .A(n36), .B(n1244), .C(n1243), .D(n33), .Z(n960) );
  COND2X1 U923 ( .A(n36), .B(n1245), .C(n1244), .D(n33), .Z(n961) );
  COND2X1 U924 ( .A(n36), .B(n1246), .C(n1245), .D(n33), .Z(n962) );
  COND2X1 U925 ( .A(n36), .B(n1247), .C(n1246), .D(n33), .Z(n963) );
  COND2X1 U926 ( .A(n36), .B(n1248), .C(n1247), .D(n33), .Z(n964) );
  COND2X1 U927 ( .A(n36), .B(n1249), .C(n1248), .D(n33), .Z(n965) );
  COND2X1 U928 ( .A(n36), .B(n1250), .C(n1249), .D(n33), .Z(n966) );
  COND2X1 U929 ( .A(n36), .B(n1251), .C(n1250), .D(n33), .Z(n967) );
  COND2X1 U930 ( .A(n36), .B(n1252), .C(n1251), .D(n33), .Z(n968) );
  COND2X1 U931 ( .A(n36), .B(n1253), .C(n1252), .D(n33), .Z(n969) );
  COND2X1 U932 ( .A(n36), .B(n1254), .C(n1253), .D(n33), .Z(n970) );
  COND2X1 U933 ( .A(n36), .B(n1255), .C(n1254), .D(n33), .Z(n971) );
  COND2X1 U934 ( .A(n36), .B(n1256), .C(n1255), .D(n33), .Z(n972) );
  COND2X1 U935 ( .A(n36), .B(n1257), .C(n1256), .D(n33), .Z(n973) );
  COND2X1 U936 ( .A(n36), .B(n1258), .C(n1257), .D(n33), .Z(n974) );
  CND2IX1 U964 ( .B(n1685), .A(n1702), .Z(n1259) );
  COND2X1 U965 ( .A(n27), .B(n1701), .C(n1288), .D(n24), .Z(n791) );
  COND2X1 U979 ( .A(n27), .B(n1274), .C(n24), .D(n1273), .Z(n989) );
  CND2IX1 U1022 ( .B(n1685), .A(n1699), .Z(n1288) );
  COND2X1 U1023 ( .A(n18), .B(n1524), .C(n1319), .D(n15), .Z(n792) );
  COND2X1 U1024 ( .A(n18), .B(n1290), .C(n15), .D(n1289), .Z(n1004) );
  COND2X1 U1025 ( .A(n18), .B(n1291), .C(n15), .D(n1290), .Z(n1005) );
  COND2X1 U1026 ( .A(n18), .B(n1292), .C(n15), .D(n1291), .Z(n1006) );
  COND2X1 U1027 ( .A(n18), .B(n1293), .C(n15), .D(n1292), .Z(n1007) );
  COND2X1 U1028 ( .A(n18), .B(n1294), .C(n15), .D(n1293), .Z(n1008) );
  COND2X1 U1029 ( .A(n18), .B(n1295), .C(n15), .D(n1294), .Z(n1009) );
  COND2X1 U1030 ( .A(n18), .B(n1296), .C(n15), .D(n1295), .Z(n1010) );
  COND2X1 U1031 ( .A(n18), .B(n1297), .C(n15), .D(n1296), .Z(n1011) );
  COND2X1 U1032 ( .A(n18), .B(n1298), .C(n15), .D(n1297), .Z(n1012) );
  COND2X1 U1033 ( .A(n18), .B(n1299), .C(n15), .D(n1298), .Z(n1013) );
  COND2X1 U1034 ( .A(n18), .B(n1300), .C(n15), .D(n1299), .Z(n1014) );
  COND2X1 U1035 ( .A(n18), .B(n1301), .C(n15), .D(n1300), .Z(n1015) );
  COND2X1 U1036 ( .A(n18), .B(n1302), .C(n15), .D(n1301), .Z(n1016) );
  COND2X1 U1037 ( .A(n18), .B(n1303), .C(n15), .D(n1302), .Z(n1017) );
  COND2X1 U1038 ( .A(n18), .B(n1304), .C(n15), .D(n1303), .Z(n1018) );
  COND2X1 U1039 ( .A(n18), .B(n1305), .C(n15), .D(n1304), .Z(n1019) );
  COND2X1 U1040 ( .A(n18), .B(n1306), .C(n15), .D(n1305), .Z(n1020) );
  COND2X1 U1041 ( .A(n18), .B(n1307), .C(n15), .D(n1306), .Z(n1021) );
  COND2X1 U1042 ( .A(n18), .B(n1308), .C(n15), .D(n1307), .Z(n1022) );
  COND2X1 U1043 ( .A(n18), .B(n1309), .C(n15), .D(n1308), .Z(n1023) );
  COND2X1 U1044 ( .A(n18), .B(n1310), .C(n15), .D(n1309), .Z(n1024) );
  COND2X1 U1045 ( .A(n18), .B(n1311), .C(n15), .D(n1310), .Z(n1025) );
  COND2X1 U1046 ( .A(n18), .B(n1312), .C(n15), .D(n1311), .Z(n1026) );
  COND2X1 U1047 ( .A(n18), .B(n1313), .C(n15), .D(n1312), .Z(n1027) );
  COND2X1 U1048 ( .A(n18), .B(n1314), .C(n15), .D(n1313), .Z(n1028) );
  COND2X1 U1049 ( .A(n18), .B(n1315), .C(n15), .D(n1314), .Z(n1029) );
  COND2X1 U1050 ( .A(n18), .B(n1316), .C(n15), .D(n1315), .Z(n1030) );
  COND2X1 U1051 ( .A(n18), .B(n1317), .C(n15), .D(n1316), .Z(n1031) );
  COND2X1 U1052 ( .A(n18), .B(n1318), .C(n15), .D(n1317), .Z(n1032) );
  CND2IX1 U1084 ( .B(n1685), .A(n1690), .Z(n1319) );
  COND2X1 U1085 ( .A(n9), .B(n1526), .C(n6), .D(n1352), .Z(n793) );
  COND2X1 U1086 ( .A(n9), .B(n1321), .C(n6), .D(n1320), .Z(n1034) );
  COND2X1 U1087 ( .A(n9), .B(n1322), .C(n6), .D(n1321), .Z(n1035) );
  COND2X1 U1088 ( .A(n9), .B(n1323), .C(n6), .D(n1322), .Z(n1036) );
  COND2X1 U1089 ( .A(n9), .B(n1324), .C(n6), .D(n1323), .Z(n1037) );
  COND2X1 U1090 ( .A(n9), .B(n1325), .C(n6), .D(n1324), .Z(n1038) );
  COND2X1 U1091 ( .A(n9), .B(n1326), .C(n6), .D(n1325), .Z(n1039) );
  COND2X1 U1092 ( .A(n9), .B(n1327), .C(n6), .D(n1326), .Z(n1040) );
  COND2X1 U1093 ( .A(n9), .B(n1328), .C(n6), .D(n1327), .Z(n1041) );
  COND2X1 U1094 ( .A(n9), .B(n1329), .C(n6), .D(n1328), .Z(n1042) );
  COND2X1 U1095 ( .A(n9), .B(n1330), .C(n6), .D(n1329), .Z(n1043) );
  COND2X1 U1096 ( .A(n9), .B(n1331), .C(n6), .D(n1330), .Z(n1044) );
  COND2X1 U1097 ( .A(n9), .B(n1332), .C(n6), .D(n1331), .Z(n1045) );
  COND2X1 U1098 ( .A(n9), .B(n1333), .C(n6), .D(n1332), .Z(n1046) );
  COND2X1 U1099 ( .A(n9), .B(n1334), .C(n6), .D(n1333), .Z(n1047) );
  COND2X1 U1100 ( .A(n9), .B(n1335), .C(n6), .D(n1334), .Z(n1048) );
  COND2X1 U1101 ( .A(n9), .B(n1336), .C(n6), .D(n1335), .Z(n1049) );
  COND2X1 U1102 ( .A(n9), .B(n1337), .C(n6), .D(n1336), .Z(n1050) );
  COND2X1 U1103 ( .A(n9), .B(n1338), .C(n6), .D(n1337), .Z(n1051) );
  COND2X1 U1104 ( .A(n9), .B(n1339), .C(n6), .D(n1338), .Z(n1052) );
  COND2X1 U1105 ( .A(n9), .B(n1340), .C(n6), .D(n1339), .Z(n1053) );
  COND2X1 U1106 ( .A(n9), .B(n1341), .C(n6), .D(n1340), .Z(n1054) );
  COND2X1 U1107 ( .A(n9), .B(n1342), .C(n6), .D(n1341), .Z(n1055) );
  COND2X1 U1108 ( .A(n9), .B(n1343), .C(n6), .D(n1342), .Z(n1056) );
  COND2X1 U1109 ( .A(n9), .B(n1344), .C(n6), .D(n1343), .Z(n1057) );
  COND2X1 U1110 ( .A(n9), .B(n1345), .C(n6), .D(n1344), .Z(n1058) );
  COND2X1 U1111 ( .A(n9), .B(n1346), .C(n6), .D(n1345), .Z(n1059) );
  COND2X1 U1112 ( .A(n9), .B(n1347), .C(n6), .D(n1346), .Z(n1060) );
  COND2X1 U1113 ( .A(n9), .B(n1348), .C(n6), .D(n1347), .Z(n1061) );
  COND2X1 U1114 ( .A(n9), .B(n1349), .C(n6), .D(n1348), .Z(n1062) );
  COND2X1 U1115 ( .A(n9), .B(n1350), .C(n6), .D(n1349), .Z(n1063) );
  COND2X1 U1116 ( .A(n9), .B(n1351), .C(n6), .D(n1350), .Z(n1064) );
  CND2IX1 U1150 ( .B(n1685), .A(n1689), .Z(n1352) );
  CENX2 U1219 ( .A(n1725), .B(a[16]), .Z(n74) );
  CENX2 U1228 ( .A(n1713), .B(a[10]), .Z(n50) );
  CFD1QXL clk_r_REG8_S1 ( .D(n348), .CP(n1679), .Q(n1670) );
  CFD1QXL clk_r_REG71_S1 ( .D(n350), .CP(n1679), .Q(n1668) );
  CFD1QXL clk_r_REG2_S1 ( .D(n347), .CP(n1679), .Q(n1671) );
  CFD1QXL clk_r_REG69_S1 ( .D(n368), .CP(n1679), .Q(n1667) );
  CFD1QXL clk_r_REG113_S1 ( .D(n278), .CP(n1679), .Q(n1677) );
  CFD1QXL clk_r_REG7_S1 ( .D(n375), .CP(n1679), .Q(n1663) );
  CFD1QXL clk_r_REG14_S1 ( .D(n399), .CP(n1679), .Q(n1659) );
  CFD1QXL clk_r_REG27_S1 ( .D(n475), .CP(n1679), .Q(n1639) );
  CFD1QXL clk_r_REG9_S1 ( .D(n426), .CP(n1679), .Q(n1653) );
  CFD1QXL clk_r_REG52_S1 ( .D(n452), .CP(n1679), .Q(n1644) );
  CFD1QXL clk_r_REG29_S1 ( .D(n499), .CP(n1679), .Q(n1634) );
  CFD1QXL clk_r_REG36_S1 ( .D(n523), .CP(n1679), .Q(n1628) );
  CFD1QXL clk_r_REG25_S1 ( .D(n503), .CP(n1679), .Q(n1630) );
  CFD1QXL clk_r_REG19_S1 ( .D(n479), .CP(n1679), .Q(n1636) );
  CFD1QXL clk_r_REG73_S1 ( .D(n620), .CP(n1679), .Q(n1600) );
  CFD1QXL clk_r_REG86_S1 ( .D(n654), .CP(n1679), .Q(n1591) );
  CFD1QXL clk_r_REG100_S1 ( .D(n721), .CP(n1679), .Q(n1568) );
  CFD1QXL clk_r_REG105_S1 ( .D(n731), .CP(n1679), .Q(n1564) );
  CFD1QXL clk_r_REG56_S1 ( .D(n584), .CP(n1679), .Q(n1610) );
  CFD1QXL clk_r_REG79_S1 ( .D(n670), .CP(n1679), .Q(n1585) );
  CFD1QXL clk_r_REG81_S1 ( .D(n656), .CP(n1679), .Q(n1589) );
  CFD1QXL clk_r_REG109_S1 ( .D(n741), .CP(n1679), .Q(n1561) );
  CFD1QXL clk_r_REG88_S1 ( .D(n684), .CP(n1679), .Q(n1582) );
  CFD1QXL clk_r_REG84_S1 ( .D(n687), .CP(n1679), .Q(n1579) );
  CFD1QXL clk_r_REG102_S1 ( .D(n722), .CP(n1679), .Q(n1567) );
  CFD1QXL clk_r_REG0_S1 ( .D(n349), .CP(n1679), .Q(n1669) );
  CFD1QXL clk_r_REG118_S1 ( .D(n287), .CP(n1679), .Q(n1674) );
  CFD1QXL clk_r_REG116_S1 ( .D(n1539), .CP(n1679), .Q(n1678) );
  CFD1QXL clk_r_REG117_S1 ( .D(n288), .CP(n1679), .Q(n1673) );
  CFD1QXL clk_r_REG13_S1 ( .D(n398), .CP(n1679), .Q(n1660) );
  CFD1QXL clk_r_REG20_S1 ( .D(n448), .CP(n1679), .Q(n1648) );
  CFD1QXL clk_r_REG39_S1 ( .D(n424), .CP(n1679), .Q(n1655) );
  CFD1QXL clk_r_REG17_S1 ( .D(n428), .CP(n1679), .Q(n1651) );
  CFD1QXL clk_r_REG18_S1 ( .D(n429), .CP(n1679), .Q(n1650) );
  CFD1QXL clk_r_REG16_S1 ( .D(n451), .CP(n1679), .Q(n1645) );
  CFD1QXL clk_r_REG22_S1 ( .D(n454), .CP(n1679), .Q(n1642) );
  CFD1QXL clk_r_REG30_S1 ( .D(n476), .CP(n1679), .Q(n1638) );
  CFD1QXL clk_r_REG55_S1 ( .D(n501), .CP(n1679), .Q(n1632) );
  CFD1QXL clk_r_REG33_S1 ( .D(n525), .CP(n1679), .Q(n1626) );
  CFD1QXL clk_r_REG32_S1 ( .D(n524), .CP(n1679), .Q(n1627) );
  CFD1QXL clk_r_REG54_S1 ( .D(n500), .CP(n1679), .Q(n1633) );
  CFD1QXL clk_r_REG59_S1 ( .D(n605), .CP(n1679), .Q(n1604) );
  CFD1QXL clk_r_REG72_S1 ( .D(n641), .CP(n1679), .Q(n1594) );
  CFD1QXL clk_r_REG49_S1 ( .D(n565), .CP(n1679), .Q(n1615) );
  CFD1QXL clk_r_REG66_S1 ( .D(n623), .CP(n1679), .Q(n1597) );
  CFD1QXL clk_r_REG57_S1 ( .D(n585), .CP(n1679), .Q(n1609) );
  CFD1QXL clk_r_REG99_S1 ( .D(n720), .CP(n1679), .Q(n1569) );
  CFD1QXL clk_r_REG110_S1 ( .D(n748), .CP(n1679), .Q(n1558) );
  CFD1QXL clk_r_REG85_S1 ( .D(n673), .CP(n1679), .Q(n1583) );
  CFD1QXL clk_r_REG90_S1 ( .D(n698), .CP(n1679), .Q(n1578) );
  CFD1QXL clk_r_REG70_S1 ( .D(n369), .CP(n1679), .Q(n1666) );
  CFD1QXL clk_r_REG4_S1 ( .D(n396), .CP(n1679), .Q(n1662) );
  CFD1QXL clk_r_REG5_S1 ( .D(n397), .CP(n1679), .Q(n1661) );
  CFD1QXL clk_r_REG11_S1 ( .D(n400), .CP(n1679), .Q(n1658) );
  CFD1QXL clk_r_REG40_S1 ( .D(n425), .CP(n1679), .Q(n1654) );
  CFD1QXL clk_r_REG28_S1 ( .D(n498), .CP(n1679), .Q(n1635) );
  CFD1QXL clk_r_REG6_S1 ( .D(n403), .CP(n1679), .Q(n1656) );
  CFD1QXL clk_r_REG96_S1 ( .D(n431), .CP(n1679), .Q(n1649) );
  CFD1QXL clk_r_REG26_S1 ( .D(n474), .CP(n1679), .Q(n1640) );
  CFD1QXL clk_r_REG23_S1 ( .D(n455), .CP(n1679), .Q(n1641) );
  CFD1QXL clk_r_REG35_S1 ( .D(n522), .CP(n1679), .Q(n1629) );
  CFD1QXL clk_r_REG41_S1 ( .D(n544), .CP(n1679), .Q(n1622) );
  CFD1QXL clk_r_REG24_S1 ( .D(n502), .CP(n1679), .Q(n1631) );
  CFD1QXL clk_r_REG37_S1 ( .D(n526), .CP(n1679), .Q(n1625) );
  CFD1QXL clk_r_REG21_S1 ( .D(n449), .CP(n1679), .Q(n1647) );
  CFD1QXL clk_r_REG87_S1 ( .D(n655), .CP(n1679), .Q(n1590) );
  CFD1QXL clk_r_REG77_S1 ( .D(n643), .CP(n1679), .Q(n1593) );
  CFD1QXL clk_r_REG89_S1 ( .D(n685), .CP(n1679), .Q(n1581) );
  CFD1QXL clk_r_REG104_S1 ( .D(n730), .CP(n1679), .Q(n1565) );
  CFD1QXL clk_r_REG91_S1 ( .D(n699), .CP(n1679), .Q(n1577) );
  CFD1QXL clk_r_REG80_S1 ( .D(n671), .CP(n1679), .Q(n1584) );
  CFD1QXL clk_r_REG101_S1 ( .D(n733), .CP(n1679), .Q(n1563) );
  CFD1QXL clk_r_REG42_S1 ( .D(n545), .CP(n1679), .Q(n1621) );
  CFD1QXL clk_r_REG44_S1 ( .D(n567), .CP(n1679), .Q(n1613) );
  CFD1QXL clk_r_REG64_S1 ( .D(n587), .CP(n1679), .Q(n1607) );
  CFD1QXL clk_r_REG122_S1 ( .D(n743), .CP(n1679), .Q(n1560) );
  CFD1QXL clk_r_REG74_S1 ( .D(n621), .CP(n1679), .Q(n1599) );
  CFD1QXL clk_r_REG112_S1 ( .D(n279), .CP(n1679), .Q(n1676) );
  CFD1QXL clk_r_REG115_S1 ( .D(n285), .CP(n1679), .Q(n1675) );
  CFD1QXL clk_r_REG120_S1 ( .D(n289), .CP(n1679), .Q(n1672) );
  CFD1QX1 clk_r_REG97_S1 ( .D(n529), .CP(n1679), .Q(n1623) );
  CFD1QX1 clk_r_REG78_S1 ( .D(n551), .CP(n1679), .Q(n1617) );
  CFD1QX2 clk_r_REG45_S1 ( .D(n546), .CP(n1679), .Q(n1620) );
  CFD1QX2 clk_r_REG34_S1 ( .D(n549), .CP(n1679), .Q(n1618) );
  CFD1QX1 clk_r_REG114_S1 ( .D(n703), .CP(n1679), .Q(n1574) );
  CFD1QX1 clk_r_REG76_S1 ( .D(n659), .CP(n1679), .Q(n1586) );
  CFD1QX1 clk_r_REG43_S1 ( .D(n566), .CP(n1679), .Q(n1614) );
  CFD1QX1 clk_r_REG46_S1 ( .D(n547), .CP(n1679), .Q(n1619) );
  CFD1QX1 clk_r_REG67_S1 ( .D(n606), .CP(n1679), .Q(n1603) );
  CFD1QX1 clk_r_REG62_S1 ( .D(n609), .CP(n1679), .Q(n1601) );
  CFD1QX1 clk_r_REG38_S1 ( .D(n527), .CP(n1679), .Q(n1624) );
  CFD1QX2 clk_r_REG83_S1 ( .D(n686), .CP(n1679), .Q(n1580) );
  CFD1QX1 clk_r_REG47_S1 ( .D(n589), .CP(n1679), .Q(n1606) );
  CFD1QX1 clk_r_REG95_S1 ( .D(n701), .CP(n1679), .Q(n1575) );
  CFD1QX1 clk_r_REG82_S1 ( .D(n657), .CP(n1679), .Q(n1588) );
  CFD1QX1 clk_r_REG50_S1 ( .D(n568), .CP(n1679), .Q(n1612) );
  CFD1QX1 clk_r_REG60_S1 ( .D(n624), .CP(n1679), .Q(n1596) );
  CFD1QXL clk_r_REG3_S1 ( .D(n371), .CP(n1679), .Q(n1665) );
  CFD1QXL clk_r_REG108_S1 ( .D(n740), .CP(n1679), .Q(n1562) );
  CFD1QXL clk_r_REG111_S1 ( .D(n746), .CP(n1679), .Q(n1559) );
  CFD1QXL clk_r_REG103_S1 ( .D(n723), .CP(n1679), .Q(n1566) );
  CFD1QXL clk_r_REG61_S1 ( .D(n625), .CP(n1679), .Q(n1595) );
  CFD1QXL clk_r_REG12_S1 ( .D(n401), .CP(n1679), .Q(n1657) );
  CFD1QXL clk_r_REG93_S1 ( .D(n711), .CP(n1679), .Q(n1572) );
  CFD1QXL clk_r_REG53_S1 ( .D(n453), .CP(n1679), .Q(n1643) );
  CFD1QXL clk_r_REG1_S1 ( .D(n373), .CP(n1679), .Q(n1664) );
  CFD1QXL clk_r_REG68_S1 ( .D(n607), .CP(n1679), .Q(n1602) );
  CFD1QXL clk_r_REG31_S1 ( .D(n477), .CP(n1679), .Q(n1637) );
  CFD1QXL clk_r_REG10_S1 ( .D(n427), .CP(n1679), .Q(n1652) );
  CFD1QXL clk_r_REG15_S1 ( .D(n450), .CP(n1679), .Q(n1646) );
  CFD1QX1 clk_r_REG107_S1 ( .D(n645), .CP(n1679), .Q(n1592) );
  CFD1QX1 clk_r_REG48_S1 ( .D(n564), .CP(n1679), .Q(n1616) );
  CFD1QX1 clk_r_REG63_S1 ( .D(n586), .CP(n1679), .Q(n1608) );
  CFD1QX1 clk_r_REG75_S1 ( .D(n658), .CP(n1679), .Q(n1587) );
  CFD1QX1 clk_r_REG98_S1 ( .D(n715), .CP(n1679), .Q(n1570) );
  CFD1QX1 clk_r_REG51_S1 ( .D(n569), .CP(n1679), .Q(n1611) );
  CFD1QX2 clk_r_REG58_S1 ( .D(n604), .CP(n1679), .Q(n1605) );
  CFD1QX1 clk_r_REG94_S1 ( .D(n700), .CP(n1679), .Q(n1576) );
  CFD1QX1 clk_r_REG106_S1 ( .D(n713), .CP(n1679), .Q(n1571) );
  CFD1QX1 clk_r_REG92_S1 ( .D(n710), .CP(n1679), .Q(n1573) );
  CFD1QX2 clk_r_REG65_S1 ( .D(n622), .CP(n1679), .Q(n1598) );
  CIVX1 U1246 ( .A(n202), .Z(n204) );
  CIVX1 U1247 ( .A(n251), .Z(n329) );
  CND2X1 U1248 ( .A(n89), .B(n1390), .Z(n91) );
  CIVX2 U1249 ( .A(a[0]), .Z(n6) );
  CNR2X1 U1250 ( .A(n579), .B(n598), .Z(n201) );
  CIVDX1 U1251 ( .A(n79), .Z0(n1522), .Z1(n1523) );
  CIVDX1 U1252 ( .A(n12), .Z0(n1524), .Z1(n1525) );
  CIVX2 U1253 ( .A(n1528), .Z(n1728) );
  CIVX1 U1254 ( .A(n1528), .Z(n1729) );
  CIVX1 U1255 ( .A(n1528), .Z(n1730) );
  CIVDX2 U1256 ( .A(n3), .Z0(n1526), .Z1(n1527) );
  CIVX2 U1257 ( .A(n1727), .Z(n1726) );
  CIVX2 U1258 ( .A(n1701), .Z(n1698) );
  CIVX2 U1259 ( .A(n1732), .Z(n1731) );
  CIVDXL U1260 ( .A(n71), .Z0(n1528), .Z1(n1529) );
  COND2XL U1261 ( .A(n27), .B(n1261), .C(n24), .D(n1260), .Z(n976) );
  COND2XL U1262 ( .A(n27), .B(n1279), .C(n24), .D(n1278), .Z(n994) );
  COND2XL U1263 ( .A(n27), .B(n1278), .C(n24), .D(n1277), .Z(n993) );
  COND2XL U1264 ( .A(n27), .B(n1282), .C(n24), .D(n1281), .Z(n997) );
  COND2XL U1265 ( .A(n27), .B(n1281), .C(n24), .D(n1280), .Z(n996) );
  COND2XL U1266 ( .A(n27), .B(n1270), .C(n24), .D(n1269), .Z(n985) );
  COND2XL U1267 ( .A(n27), .B(n1269), .C(n24), .D(n1268), .Z(n984) );
  COND2XL U1268 ( .A(n27), .B(n1264), .C(n24), .D(n1263), .Z(n979) );
  COND2XL U1269 ( .A(n27), .B(n1266), .C(n24), .D(n1265), .Z(n981) );
  COND2XL U1270 ( .A(n27), .B(n1273), .C(n24), .D(n1272), .Z(n988) );
  COND2XL U1271 ( .A(n27), .B(n1272), .C(n24), .D(n1271), .Z(n987) );
  COND2XL U1272 ( .A(n27), .B(n1262), .C(n24), .D(n1261), .Z(n977) );
  COND2XL U1273 ( .A(n27), .B(n1265), .C(n24), .D(n1264), .Z(n980) );
  COND2XL U1274 ( .A(n27), .B(n1271), .C(n24), .D(n1270), .Z(n986) );
  COND2XL U1275 ( .A(n27), .B(n1268), .C(n24), .D(n1267), .Z(n983) );
  COND2XL U1276 ( .A(n27), .B(n1286), .C(n24), .D(n1285), .Z(n1001) );
  COND2XL U1277 ( .A(n27), .B(n1280), .C(n24), .D(n1279), .Z(n995) );
  COND2XL U1278 ( .A(n27), .B(n1276), .C(n24), .D(n1275), .Z(n991) );
  COND2XL U1279 ( .A(n27), .B(n1285), .C(n24), .D(n1284), .Z(n1000) );
  COND2XL U1280 ( .A(n27), .B(n1277), .C(n24), .D(n1276), .Z(n992) );
  COND2XL U1281 ( .A(n27), .B(n1263), .C(n24), .D(n1262), .Z(n978) );
  COND2XL U1282 ( .A(n27), .B(n1283), .C(n24), .D(n1282), .Z(n998) );
  COND2XL U1283 ( .A(n27), .B(n1275), .C(n24), .D(n1274), .Z(n990) );
  COND2XL U1284 ( .A(n27), .B(n1267), .C(n24), .D(n1266), .Z(n982) );
  COND2XL U1285 ( .A(n27), .B(n1284), .C(n24), .D(n1283), .Z(n999) );
  COND2X1 U1286 ( .A(n27), .B(n1287), .C(n24), .D(n1286), .Z(n1002) );
  CND2X2 U1287 ( .A(n1396), .B(n42), .Z(n44) );
  CHA1XL U1288 ( .A(n789), .B(n1026), .CO(n752), .S(n753) );
  CFA1XL U1289 ( .A(n823), .B(n845), .CI(n833), .CO(n576), .S(n577) );
  COND2XL U1290 ( .A(n91), .B(n1101), .C(n1100), .D(n89), .Z(n824) );
  COND2XL U1291 ( .A(n91), .B(n1103), .C(n1102), .D(n89), .Z(n826) );
  COND2XL U1292 ( .A(n91), .B(n1105), .C(n1104), .D(n89), .Z(n828) );
  COND2XL U1293 ( .A(n91), .B(n1104), .C(n1103), .D(n89), .Z(n827) );
  COND2XL U1294 ( .A(n91), .B(n1106), .C(n1105), .D(n89), .Z(n829) );
  COND2XL U1295 ( .A(n1111), .B(n91), .C(n1110), .D(n89), .Z(n834) );
  COND2XL U1296 ( .A(n91), .B(n1109), .C(n1108), .D(n89), .Z(n832) );
  COND2XL U1297 ( .A(n91), .B(n1102), .C(n1101), .D(n89), .Z(n825) );
  COND2XL U1298 ( .A(n91), .B(n1736), .C(n89), .D(n1112), .Z(n783) );
  COND2XL U1299 ( .A(n91), .B(n1107), .C(n1106), .D(n89), .Z(n830) );
  CND2X4 U1300 ( .A(n1392), .B(n74), .Z(n77) );
  CEOX1 U1301 ( .A(a[16]), .B(n1529), .Z(n1392) );
  CANR1X1 U1302 ( .A(n175), .B(n1544), .C(n170), .Z(n168) );
  CENXL U1303 ( .A(n1697), .B(b[27]), .Z(n1260) );
  COND2XL U1304 ( .A(n69), .B(n1146), .C(n1145), .D(n66), .Z(n866) );
  COND2XL U1305 ( .A(n69), .B(n1158), .C(n1157), .D(n66), .Z(n878) );
  COND2XL U1306 ( .A(n69), .B(n1727), .C(n1163), .D(n66), .Z(n786) );
  COND2XL U1307 ( .A(n69), .B(n1149), .C(n1148), .D(n66), .Z(n869) );
  COND2XL U1308 ( .A(n69), .B(n1156), .C(n1155), .D(n66), .Z(n876) );
  COND2XL U1309 ( .A(n69), .B(n1154), .C(n1153), .D(n66), .Z(n874) );
  COND2XL U1310 ( .A(n69), .B(n1150), .C(n1149), .D(n66), .Z(n870) );
  COND2XL U1311 ( .A(n69), .B(n1151), .C(n1150), .D(n66), .Z(n871) );
  COND2XL U1312 ( .A(n69), .B(n1157), .C(n1156), .D(n66), .Z(n877) );
  CENXL U1313 ( .A(n1722), .B(n1373), .Z(n1172) );
  CENX2 U1314 ( .A(n1722), .B(a[14]), .Z(n66) );
  COND1X2 U1315 ( .A(n195), .B(n182), .C(n183), .Z(n181) );
  CANR1X2 U1316 ( .A(n204), .B(n1542), .C(n197), .Z(n195) );
  CIVXL U1317 ( .A(n208), .Z(n207) );
  CENXL U1318 ( .A(n1695), .B(b[26]), .Z(n1261) );
  COND1X1 U1319 ( .A(n209), .B(n221), .C(n210), .Z(n208) );
  CANR1X1 U1320 ( .A(n241), .B(n222), .C(n223), .Z(n221) );
  CIVXL U1321 ( .A(n241), .Z(n240) );
  CIVDX1 U1322 ( .A(n1742), .Z1(product[7]) );
  CEOX1 U1323 ( .A(n1726), .B(a[14]), .Z(n1537) );
  CENXL U1324 ( .A(n1534), .B(n121), .Z(product[29]) );
  CANR1X1 U1325 ( .A(n237), .B(n1552), .C(n230), .Z(n228) );
  CENXL U1326 ( .A(n1722), .B(n1374), .Z(n1173) );
  CENXL U1327 ( .A(n1726), .B(n1374), .Z(n1152) );
  CENXL U1328 ( .A(n1729), .B(n1374), .Z(n1133) );
  CENXL U1329 ( .A(n1731), .B(n1374), .Z(n1116) );
  CENXL U1330 ( .A(n1698), .B(n1374), .Z(n1277) );
  CENXL U1331 ( .A(n1527), .B(n1374), .Z(n1341) );
  CENXL U1332 ( .A(n1694), .B(n1374), .Z(n1308) );
  CENXL U1333 ( .A(n1715), .B(n1374), .Z(n1221) );
  CENXL U1334 ( .A(n1734), .B(n1374), .Z(n1101) );
  CENXL U1335 ( .A(n1706), .B(n1374), .Z(n1248) );
  CEOX2 U1336 ( .A(a[6]), .B(n1707), .Z(n1397) );
  CANR1XL U1337 ( .A(n1545), .B(n158), .C(n155), .Z(n1531) );
  CANR1XL U1338 ( .A(n1546), .B(n1533), .C(n163), .Z(n1532) );
  COND1X1 U1339 ( .A(n159), .B(n161), .C(n160), .Z(n158) );
  CANR1X1 U1340 ( .A(n1545), .B(n158), .C(n155), .Z(n153) );
  CANR1X1 U1341 ( .A(n1546), .B(n1533), .C(n163), .Z(n161) );
  CIVX1 U1342 ( .A(n199), .Z(n197) );
  CIVX1 U1343 ( .A(n201), .Z(n322) );
  COND1XL U1344 ( .A(n167), .B(n179), .C(n168), .Z(n166) );
  CENXL U1345 ( .A(n1688), .B(b[25]), .Z(n1326) );
  CENXL U1346 ( .A(n1700), .B(b[25]), .Z(n1262) );
  CENXL U1347 ( .A(n1694), .B(b[25]), .Z(n1293) );
  CANR1X2 U1348 ( .A(n190), .B(n1543), .C(n185), .Z(n183) );
  CANR1X1 U1349 ( .A(n217), .B(n1553), .C(n212), .Z(n210) );
  CENXL U1350 ( .A(n1536), .B(n150), .Z(product[31]) );
  CENXL U1351 ( .A(n1688), .B(b[24]), .Z(n1327) );
  CENXL U1352 ( .A(n1695), .B(b[24]), .Z(n1263) );
  CENXL U1353 ( .A(n1694), .B(b[24]), .Z(n1294) );
  CENXL U1354 ( .A(n1702), .B(b[24]), .Z(n1234) );
  CANR1X2 U1355 ( .A(n180), .B(n208), .C(n181), .Z(n179) );
  CNR2X1 U1356 ( .A(n182), .B(n194), .Z(n180) );
  CIVX1 U1357 ( .A(n21), .Z(n1701) );
  CEOX2 U1358 ( .A(n1698), .B(a[6]), .Z(n1554) );
  CIVX4 U1359 ( .A(n1554), .Z(n33) );
  COND1X1 U1360 ( .A(n167), .B(n179), .C(n168), .Z(n1533) );
  CANR1X1 U1361 ( .A(n260), .B(n268), .C(n261), .Z(n259) );
  COND1X1 U1362 ( .A(n257), .B(n251), .C(n252), .Z(n250) );
  COND2X1 U1363 ( .A(n84), .B(n1125), .C(n1124), .D(n82), .Z(n847) );
  CEOX2 U1364 ( .A(n1705), .B(a[8]), .Z(n1557) );
  CIVX2 U1365 ( .A(n1709), .Z(n1705) );
  CENXL U1366 ( .A(n1705), .B(n1376), .Z(n1250) );
  COND2XL U1367 ( .A(n44), .B(n1718), .C(n1232), .D(n42), .Z(n789) );
  COND2X1 U1368 ( .A(n44), .B(n1230), .C(n1229), .D(n42), .Z(n947) );
  CENXL U1369 ( .A(n1705), .B(b[25]), .Z(n1233) );
  COND2XL U1370 ( .A(n44), .B(n1223), .C(n1222), .D(n42), .Z(n940) );
  CIVX1 U1371 ( .A(n1727), .Z(n1725) );
  CENXL U1372 ( .A(n1725), .B(n1378), .Z(n1156) );
  CND2IXL U1373 ( .B(n1685), .A(n1725), .Z(n1163) );
  CIVXL U1374 ( .A(n179), .Z(n178) );
  CEOX1 U1375 ( .A(a[10]), .B(n1720), .Z(n1395) );
  CIVX1 U1376 ( .A(n1721), .Z(n1720) );
  CENXL U1377 ( .A(n1720), .B(n1366), .Z(n1188) );
  CENXL U1378 ( .A(n1720), .B(n1369), .Z(n1191) );
  CENXL U1379 ( .A(n1720), .B(n1368), .Z(n1190) );
  CENXL U1380 ( .A(n1720), .B(n1373), .Z(n1195) );
  CENXL U1381 ( .A(n1720), .B(n1370), .Z(n1192) );
  CENXL U1382 ( .A(n1720), .B(n1374), .Z(n1196) );
  CENXL U1383 ( .A(n1720), .B(n1367), .Z(n1189) );
  COND1X1 U1384 ( .A(n259), .B(n242), .C(n243), .Z(n241) );
  CND2XL U1385 ( .A(n249), .B(n1551), .Z(n242) );
  CANR1X1 U1386 ( .A(n1551), .B(n250), .C(n245), .Z(n243) );
  COND1X1 U1387 ( .A(n151), .B(n153), .C(n152), .Z(n150) );
  CEOX1 U1388 ( .A(a[2]), .B(n1525), .Z(n1399) );
  CIVX4 U1389 ( .A(n1526), .Z(n1689) );
  CIVX1 U1390 ( .A(n1526), .Z(n1688) );
  COND2XL U1391 ( .A(n53), .B(n1203), .C(n1202), .D(n50), .Z(n921) );
  CENX4 U1392 ( .A(n1719), .B(a[12]), .Z(n58) );
  CNR2XL U1393 ( .A(n224), .B(n227), .Z(n222) );
  CIVX1 U1394 ( .A(n1724), .Z(n1723) );
  CIVX2 U1395 ( .A(n1739), .Z(n1738) );
  CNR2XL U1396 ( .A(n251), .B(n256), .Z(n249) );
  COND2XL U1397 ( .A(n69), .B(n1161), .C(n1160), .D(n66), .Z(n881) );
  CND2X4 U1398 ( .A(n1394), .B(n58), .Z(n61) );
  CEOX2 U1399 ( .A(a[12]), .B(n1723), .Z(n1394) );
  COND1XL U1400 ( .A(n159), .B(n1532), .C(n160), .Z(n1534) );
  CAOR1XL U1401 ( .A(n241), .B(n222), .C(n223), .Z(n1535) );
  CND2X1 U1402 ( .A(n1543), .B(n1540), .Z(n182) );
  CANR1XL U1403 ( .A(n302), .B(n1548), .C(n299), .Z(n297) );
  CANR1XL U1404 ( .A(n310), .B(n1549), .C(n307), .Z(n305) );
  CND2X2 U1405 ( .A(n1537), .B(n66), .Z(n69) );
  CEOXL U1406 ( .A(n1531), .B(n120), .Z(product[30]) );
  CEOXL U1407 ( .A(n124), .B(n173), .Z(product[26]) );
  CND2XL U1408 ( .A(n1544), .B(n172), .Z(n124) );
  CEOXL U1409 ( .A(n126), .B(n188), .Z(product[24]) );
  CND2XL U1410 ( .A(n1543), .B(n187), .Z(n126) );
  CND2XL U1411 ( .A(n315), .B(n160), .Z(n122) );
  CND2XL U1412 ( .A(n322), .B(n202), .Z(n129) );
  CEOXL U1413 ( .A(n297), .B(n145), .Z(product[5]) );
  CND2XL U1414 ( .A(n1548), .B(n301), .Z(n146) );
  CND2XL U1415 ( .A(n1549), .B(n309), .Z(n148) );
  CND2XL U1416 ( .A(n1545), .B(n157), .Z(n121) );
  CND2XL U1417 ( .A(n1546), .B(n165), .Z(n123) );
  CND2XL U1418 ( .A(n1541), .B(n177), .Z(n125) );
  CND2XL U1419 ( .A(n1540), .B(n192), .Z(n127) );
  CND2XL U1420 ( .A(n1542), .B(n322), .Z(n194) );
  CNR2XL U1421 ( .A(n747), .B(n754), .Z(n278) );
  CND2XL U1422 ( .A(n755), .B(n760), .Z(n285) );
  CNR2XL U1423 ( .A(n262), .B(n265), .Z(n260) );
  CEOXL U1424 ( .A(n130), .B(n215), .Z(product[20]) );
  CND2XL U1425 ( .A(n1553), .B(n214), .Z(n130) );
  CND2XL U1426 ( .A(n332), .B(n266), .Z(n139) );
  CND2XL U1427 ( .A(n1551), .B(n247), .Z(n135) );
  CND2XL U1428 ( .A(n327), .B(n235), .Z(n134) );
  CND2XL U1429 ( .A(n330), .B(n257), .Z(n137) );
  CND2XL U1430 ( .A(n1552), .B(n232), .Z(n133) );
  CND2XL U1431 ( .A(n325), .B(n225), .Z(n132) );
  CND2XL U1432 ( .A(n1550), .B(n219), .Z(n131) );
  CND2XL U1433 ( .A(n777), .B(n792), .Z(n304) );
  CND2XL U1434 ( .A(n1552), .B(n327), .Z(n227) );
  CNR2XL U1435 ( .A(n761), .B(n766), .Z(n287) );
  COR2XL U1436 ( .A(n1063), .B(n1033), .Z(n1549) );
  CND2IXL U1437 ( .B(n311), .A(n312), .Z(n149) );
  CENX1 U1438 ( .A(n343), .B(n358), .Z(n1536) );
  CND2XL U1439 ( .A(n695), .B(n706), .Z(n252) );
  CND2XL U1440 ( .A(n1555), .B(n274), .Z(n140) );
  CNR2IXL U1441 ( .B(n1685), .A(n95), .Z(n823) );
  COND2XL U1442 ( .A(n91), .B(n1110), .C(n1109), .D(n89), .Z(n833) );
  CNR2IXL U1443 ( .B(n1685), .A(n110), .Z(n799) );
  COND2XL U1444 ( .A(n1077), .B(n107), .C(n105), .D(n1076), .Z(n803) );
  CNR2IXL U1445 ( .B(n1685), .A(n42), .Z(n949) );
  CNR2IXL U1446 ( .B(n1685), .A(n89), .Z(n835) );
  CNR2IXL U1447 ( .B(n1685), .A(n66), .Z(n883) );
  CNR2IXL U1448 ( .B(n1685), .A(n100), .Z(n813) );
  COND2XL U1449 ( .A(n91), .B(n1108), .C(n1107), .D(n89), .Z(n831) );
  CND2XL U1450 ( .A(n719), .B(n728), .Z(n263) );
  CNR2IXL U1451 ( .B(n1685), .A(n6), .Z(product[0]) );
  COND2XL U1452 ( .A(n102), .B(n1081), .C(n100), .D(n1080), .Z(n806) );
  COND2XL U1453 ( .A(n53), .B(n1200), .C(n1199), .D(n50), .Z(n918) );
  CENX2 U1454 ( .A(n1728), .B(a[18]), .Z(n82) );
  CND2IX4 U1455 ( .B(n1538), .A(n6), .Z(n9) );
  CENXL U1456 ( .A(a[0]), .B(n1689), .Z(n1538) );
  CND2X2 U1457 ( .A(n1391), .B(n82), .Z(n84) );
  CNIVX1 U1458 ( .A(n1382), .Z(n1680) );
  CNIVX1 U1459 ( .A(n1381), .Z(n1681) );
  CNIVX1 U1460 ( .A(n1379), .Z(n1683) );
  CNIVX1 U1461 ( .A(n1380), .Z(n1682) );
  CIVX3 U1462 ( .A(n1556), .Z(n24) );
  CEOXL U1463 ( .A(a[8]), .B(n1716), .Z(n1396) );
  CND2X2 U1464 ( .A(n95), .B(n1389), .Z(n97) );
  COND2XL U1465 ( .A(n1067), .B(n114), .C(n1410), .D(n115), .Z(n778) );
  CND2IXL U1466 ( .B(n1685), .A(n113), .Z(n1067) );
  CIVX3 U1467 ( .A(n1557), .Z(n42) );
  CNIVXL U1468 ( .A(n1383), .Z(n1687) );
  CND2XL U1469 ( .A(n1385), .B(n114), .Z(n115) );
  CND2IXL U1470 ( .B(n1685), .A(n109), .Z(n1072) );
  COND1XL U1471 ( .A(n194), .B(n207), .C(n195), .Z(n193) );
  CND2X1 U1472 ( .A(n1544), .B(n1541), .Z(n167) );
  COND1XL U1473 ( .A(n297), .B(n295), .C(n296), .Z(n294) );
  COND1XL U1474 ( .A(n305), .B(n303), .C(n304), .Z(n302) );
  CENX1 U1475 ( .A(n200), .B(n128), .Z(product[22]) );
  CND2X1 U1476 ( .A(n1542), .B(n199), .Z(n128) );
  COND1XL U1477 ( .A(n201), .B(n207), .C(n202), .Z(n200) );
  CANR1XL U1478 ( .A(n294), .B(n1547), .C(n291), .Z(n289) );
  CENX1 U1479 ( .A(n144), .B(n294), .Z(product[6]) );
  CND2X1 U1480 ( .A(n1547), .B(n293), .Z(n144) );
  CENX1 U1481 ( .A(n146), .B(n302), .Z(product[4]) );
  CENX1 U1482 ( .A(n148), .B(n310), .Z(product[2]) );
  CENX1 U1483 ( .A(n193), .B(n127), .Z(product[23]) );
  CENX1 U1484 ( .A(n178), .B(n125), .Z(product[25]) );
  CENX1 U1485 ( .A(n166), .B(n123), .Z(product[27]) );
  CND2X1 U1486 ( .A(n338), .B(n296), .Z(n145) );
  CEOXL U1487 ( .A(n305), .B(n147), .Z(product[3]) );
  CND2X1 U1488 ( .A(n340), .B(n304), .Z(n147) );
  CND2X1 U1489 ( .A(n313), .B(n152), .Z(n120) );
  CEOXL U1490 ( .A(n122), .B(n1532), .Z(product[28]) );
  CANR1XL U1491 ( .A(n1541), .B(n178), .C(n175), .Z(n173) );
  CANR1XL U1492 ( .A(n1540), .B(n193), .C(n190), .Z(n188) );
  CEOXL U1493 ( .A(n129), .B(n207), .Z(product[21]) );
  CND2XL U1494 ( .A(n747), .B(n754), .Z(n279) );
  COR2X1 U1495 ( .A(n755), .B(n760), .Z(n1539) );
  CANR1XL U1496 ( .A(n1550), .B(n1535), .C(n217), .Z(n215) );
  CEOX1 U1497 ( .A(n135), .B(n248), .Z(product[15]) );
  CANR1XL U1498 ( .A(n249), .B(n258), .C(n250), .Z(n248) );
  COND1XL U1499 ( .A(n266), .B(n262), .C(n263), .Z(n261) );
  COND1XL U1500 ( .A(n228), .B(n224), .C(n225), .Z(n223) );
  CND2X1 U1501 ( .A(n1553), .B(n1550), .Z(n209) );
  CENX1 U1502 ( .A(n264), .B(n138), .Z(product[12]) );
  CND2X1 U1503 ( .A(n331), .B(n263), .Z(n138) );
  COND1XL U1504 ( .A(n265), .B(n267), .C(n266), .Z(n264) );
  CENX1 U1505 ( .A(n258), .B(n137), .Z(product[13]) );
  CENX1 U1506 ( .A(n233), .B(n133), .Z(product[17]) );
  COND1XL U1507 ( .A(n234), .B(n240), .C(n235), .Z(n233) );
  CENX1 U1508 ( .A(n226), .B(n132), .Z(product[18]) );
  COND1XL U1509 ( .A(n227), .B(n240), .C(n228), .Z(n226) );
  CENX1 U1510 ( .A(n1535), .B(n131), .Z(product[19]) );
  CNR2X1 U1511 ( .A(n415), .B(n440), .Z(n159) );
  CNR2X1 U1512 ( .A(n359), .B(n386), .Z(n151) );
  CNR2X1 U1513 ( .A(n771), .B(n774), .Z(n295) );
  CNR2X1 U1514 ( .A(n777), .B(n792), .Z(n303) );
  CEOX1 U1515 ( .A(n139), .B(n267), .Z(product[11]) );
  CEOX1 U1516 ( .A(n136), .B(n253), .Z(product[14]) );
  CND2X1 U1517 ( .A(n329), .B(n252), .Z(n136) );
  CANR1XL U1518 ( .A(n330), .B(n258), .C(n255), .Z(n253) );
  CEOX1 U1519 ( .A(n134), .B(n240), .Z(product[16]) );
  COR2X1 U1520 ( .A(n537), .B(n558), .Z(n1540) );
  COR2X1 U1521 ( .A(n491), .B(n514), .Z(n1541) );
  COR2X1 U1522 ( .A(n559), .B(n578), .Z(n1542) );
  CND2X1 U1523 ( .A(n579), .B(n598), .Z(n202) );
  COR2X1 U1524 ( .A(n515), .B(n536), .Z(n1543) );
  COR2X1 U1525 ( .A(n467), .B(n490), .Z(n1544) );
  CND2X1 U1526 ( .A(n537), .B(n558), .Z(n192) );
  CND2X1 U1527 ( .A(n515), .B(n536), .Z(n187) );
  CND2X1 U1528 ( .A(n559), .B(n578), .Z(n199) );
  CND2X1 U1529 ( .A(n491), .B(n514), .Z(n177) );
  CND2X1 U1530 ( .A(n467), .B(n490), .Z(n172) );
  CND2X1 U1531 ( .A(n775), .B(n776), .Z(n301) );
  CND2X1 U1532 ( .A(n767), .B(n770), .Z(n293) );
  CND2X1 U1533 ( .A(n387), .B(n414), .Z(n157) );
  CND2X1 U1534 ( .A(n441), .B(n466), .Z(n165) );
  CND2X1 U1535 ( .A(n1064), .B(n793), .Z(n312) );
  CND2X1 U1536 ( .A(n1063), .B(n1033), .Z(n309) );
  CND2X1 U1537 ( .A(n771), .B(n774), .Z(n296) );
  CND2X1 U1538 ( .A(n415), .B(n440), .Z(n160) );
  CND2X1 U1539 ( .A(n359), .B(n386), .Z(n152) );
  COR2X1 U1540 ( .A(n387), .B(n414), .Z(n1545) );
  COR2X1 U1541 ( .A(n441), .B(n466), .Z(n1546) );
  COR2X1 U1542 ( .A(n767), .B(n770), .Z(n1547) );
  COR2X1 U1543 ( .A(n775), .B(n776), .Z(n1548) );
  CND2XL U1544 ( .A(n761), .B(n766), .Z(n288) );
  CNR2XL U1545 ( .A(n1064), .B(n793), .Z(n311) );
  CENX1 U1546 ( .A(n1684), .B(n1689), .Z(n1351) );
  CNR2IX1 U1547 ( .B(n1685), .A(n114), .Z(n795) );
  CIVX2 U1548 ( .A(n1741), .Z(n1740) );
  COND1XL U1549 ( .A(n281), .B(n269), .C(n270), .Z(n268) );
  CND2X1 U1550 ( .A(n1555), .B(n334), .Z(n269) );
  CANR1XL U1551 ( .A(n277), .B(n1555), .C(n272), .Z(n270) );
  CNR2X1 U1552 ( .A(n729), .B(n738), .Z(n265) );
  CIVX2 U1553 ( .A(n1721), .Z(n1719) );
  CNR2X1 U1554 ( .A(n695), .B(n706), .Z(n251) );
  CNR2X1 U1555 ( .A(n635), .B(n650), .Z(n224) );
  CNR2X1 U1556 ( .A(n719), .B(n728), .Z(n262) );
  CNR2IXL U1557 ( .B(n1685), .A(n15), .Z(n1033) );
  CENX1 U1558 ( .A(n1726), .B(n1686), .Z(n1161) );
  CENX1 U1559 ( .A(n1726), .B(n1680), .Z(n1160) );
  CENX1 U1560 ( .A(n1726), .B(n1681), .Z(n1159) );
  CENX1 U1561 ( .A(n1731), .B(n1686), .Z(n1125) );
  CENX1 U1562 ( .A(n1728), .B(n1681), .Z(n1140) );
  CENX1 U1563 ( .A(n1725), .B(n1683), .Z(n1157) );
  CENX1 U1564 ( .A(n1728), .B(n1682), .Z(n1139) );
  CENX1 U1565 ( .A(n1731), .B(n1680), .Z(n1124) );
  CENX1 U1566 ( .A(n1728), .B(n1683), .Z(n1138) );
  CENX1 U1567 ( .A(n1686), .B(n1735), .Z(n1110) );
  CENX1 U1568 ( .A(n1731), .B(n1681), .Z(n1123) );
  CENX1 U1569 ( .A(n1523), .B(n1682), .Z(n1122) );
  CENX1 U1570 ( .A(n1680), .B(n1735), .Z(n1109) );
  CENX1 U1571 ( .A(n1523), .B(n1683), .Z(n1121) );
  CENX1 U1572 ( .A(n1681), .B(n1735), .Z(n1108) );
  CENX1 U1573 ( .A(n1704), .B(n1681), .Z(n1255) );
  CENX1 U1574 ( .A(n1713), .B(n1680), .Z(n1229) );
  CENX1 U1575 ( .A(n1713), .B(n1681), .Z(n1228) );
  CENX1 U1576 ( .A(n1704), .B(n1683), .Z(n1253) );
  CENX1 U1577 ( .A(n1704), .B(n1682), .Z(n1254) );
  CENX1 U1578 ( .A(n1729), .B(n1686), .Z(n1142) );
  CENX1 U1579 ( .A(n1704), .B(n1680), .Z(n1256) );
  CENX1 U1580 ( .A(n1705), .B(n1686), .Z(n1257) );
  CENX1 U1581 ( .A(n1725), .B(n1682), .Z(n1158) );
  CENX1 U1582 ( .A(n1728), .B(n1680), .Z(n1141) );
  CENX1 U1583 ( .A(n1713), .B(n1686), .Z(n1230) );
  CENX1 U1584 ( .A(n1719), .B(n1686), .Z(n1205) );
  CENX1 U1585 ( .A(n1719), .B(n1682), .Z(n1202) );
  CENX1 U1586 ( .A(n1722), .B(n1680), .Z(n1181) );
  CENX1 U1587 ( .A(n1722), .B(n1681), .Z(n1180) );
  CENX1 U1588 ( .A(n1722), .B(n1682), .Z(n1179) );
  CENX1 U1589 ( .A(n1722), .B(n1683), .Z(n1178) );
  CENX1 U1590 ( .A(n1682), .B(n1735), .Z(n1107) );
  CENX1 U1591 ( .A(n1683), .B(n1735), .Z(n1106) );
  CENX1 U1592 ( .A(n1722), .B(n1686), .Z(n1182) );
  CENX1 U1593 ( .A(n1719), .B(n1680), .Z(n1204) );
  CENX1 U1594 ( .A(n1719), .B(n1681), .Z(n1203) );
  CENX1 U1595 ( .A(n1712), .B(n1682), .Z(n1227) );
  CENX1 U1596 ( .A(n1712), .B(n1683), .Z(n1226) );
  CENX1 U1597 ( .A(n1719), .B(n1683), .Z(n1201) );
  CENX1 U1598 ( .A(n1527), .B(n1680), .Z(n1349) );
  CENX1 U1599 ( .A(n1527), .B(n1681), .Z(n1348) );
  CENX1 U1600 ( .A(n1527), .B(n1682), .Z(n1347) );
  CENX1 U1601 ( .A(n1697), .B(n1687), .Z(n1286) );
  CENX1 U1602 ( .A(n1527), .B(n1683), .Z(n1346) );
  CENX1 U1603 ( .A(n1696), .B(n1682), .Z(n1283) );
  CENX1 U1604 ( .A(n1683), .B(n1740), .Z(n1082) );
  CENX1 U1605 ( .A(n1697), .B(n1680), .Z(n1285) );
  CENX1 U1606 ( .A(n1692), .B(n1681), .Z(n1315) );
  CENX1 U1607 ( .A(n1692), .B(n1682), .Z(n1314) );
  CENX1 U1608 ( .A(n1692), .B(n1680), .Z(n1316) );
  CENX1 U1609 ( .A(n1692), .B(n1683), .Z(n1313) );
  CENX1 U1610 ( .A(n1527), .B(n1687), .Z(n1350) );
  CENX1 U1611 ( .A(n1697), .B(n1681), .Z(n1284) );
  CENX1 U1612 ( .A(n1693), .B(n1687), .Z(n1317) );
  CENX1 U1613 ( .A(n1680), .B(n1738), .Z(n1096) );
  CENX1 U1614 ( .A(n1686), .B(n1738), .Z(n1097) );
  CENX1 U1615 ( .A(n1681), .B(n1738), .Z(n1095) );
  CENX1 U1616 ( .A(n1686), .B(n1740), .Z(n1086) );
  CENX1 U1617 ( .A(n1682), .B(n1738), .Z(n1094) );
  CENX1 U1618 ( .A(n1680), .B(n1740), .Z(n1085) );
  CENX1 U1619 ( .A(n1683), .B(n1738), .Z(n1093) );
  CENX1 U1620 ( .A(n1681), .B(n1740), .Z(n1084) );
  CENX1 U1621 ( .A(n1682), .B(n1740), .Z(n1083) );
  CENX1 U1622 ( .A(n1696), .B(n1683), .Z(n1282) );
  CNR2X1 U1623 ( .A(n707), .B(n718), .Z(n256) );
  CIVX2 U1624 ( .A(n1724), .Z(n1722) );
  CENX1 U1625 ( .A(n1684), .B(n1707), .Z(n1258) );
  CENX1 U1626 ( .A(n1684), .B(n1726), .Z(n1162) );
  CENX1 U1627 ( .A(n1684), .B(n1716), .Z(n1231) );
  CENX1 U1628 ( .A(n1684), .B(n1720), .Z(n1206) );
  CENX1 U1629 ( .A(n1685), .B(n1723), .Z(n1183) );
  CENX1 U1630 ( .A(n1684), .B(n1735), .Z(n1111) );
  CENX1 U1631 ( .A(n1684), .B(n1731), .Z(n1126) );
  CENX1 U1632 ( .A(n1684), .B(n1738), .Z(n1098) );
  CENX1 U1633 ( .A(n1684), .B(n1740), .Z(n1087) );
  CNR2IX1 U1634 ( .B(n1685), .A(n24), .Z(n1003) );
  CENX1 U1635 ( .A(n1685), .B(n1700), .Z(n1287) );
  CENX1 U1636 ( .A(n1684), .B(n1525), .Z(n1318) );
  CNR2X1 U1637 ( .A(n667), .B(n680), .Z(n234) );
  CNR2IX1 U1638 ( .B(n1685), .A(n58), .Z(n903) );
  CNR2IXL U1639 ( .B(n1685), .A(n74), .Z(n865) );
  CNR2IX1 U1640 ( .B(n1685), .A(n82), .Z(n849) );
  COR2X1 U1641 ( .A(n617), .B(n634), .Z(n1550) );
  COR2X1 U1642 ( .A(n681), .B(n694), .Z(n1551) );
  COR2X1 U1643 ( .A(n651), .B(n666), .Z(n1552) );
  CND2X1 U1644 ( .A(n667), .B(n680), .Z(n235) );
  COR2X1 U1645 ( .A(n599), .B(n616), .Z(n1553) );
  CND2X1 U1646 ( .A(n707), .B(n718), .Z(n257) );
  CNR2IXL U1647 ( .B(n1685), .A(n50), .Z(n925) );
  CNR2IX1 U1648 ( .B(n1685), .A(n33), .Z(n975) );
  CNR2IX1 U1649 ( .B(n1685), .A(n105), .Z(n805) );
  CND2X1 U1650 ( .A(n729), .B(n738), .Z(n266) );
  CND2X1 U1651 ( .A(n617), .B(n634), .Z(n219) );
  CND2X1 U1652 ( .A(n651), .B(n666), .Z(n232) );
  CND2X1 U1653 ( .A(n681), .B(n694), .Z(n247) );
  CND2X1 U1654 ( .A(n599), .B(n616), .Z(n214) );
  CEOX1 U1655 ( .A(n806), .B(n796), .Z(n357) );
  CND2X1 U1656 ( .A(n635), .B(n650), .Z(n225) );
  CENX1 U1657 ( .A(n1685), .B(n1529), .Z(n1143) );
  CEOX1 U1658 ( .A(n275), .B(n140), .Z(product[10]) );
  CANR1XL U1659 ( .A(n334), .B(n280), .C(n277), .Z(n275) );
  CENX1 U1660 ( .A(n1523), .B(a[20]), .Z(n89) );
  CENX1 U1661 ( .A(n1733), .B(a[22]), .Z(n95) );
  CENX1 U1662 ( .A(n1738), .B(a[24]), .Z(n100) );
  CENX1 U1663 ( .A(n1740), .B(a[26]), .Z(n105) );
  CENX1 U1664 ( .A(n1712), .B(n1377), .Z(n1224) );
  CENX1 U1665 ( .A(n1722), .B(n1378), .Z(n1177) );
  CENX1 U1666 ( .A(n1726), .B(n1376), .Z(n1154) );
  CENX1 U1667 ( .A(n1731), .B(n1372), .Z(n1114) );
  CENX1 U1668 ( .A(n1712), .B(n1378), .Z(n1225) );
  CENX1 U1669 ( .A(n1728), .B(n1378), .Z(n1137) );
  CENX1 U1670 ( .A(n1523), .B(n1378), .Z(n1120) );
  CENX1 U1671 ( .A(n1730), .B(n1376), .Z(n1135) );
  CENX1 U1672 ( .A(n1731), .B(n1377), .Z(n1119) );
  CENX1 U1673 ( .A(n1714), .B(n1376), .Z(n1223) );
  CENX1 U1674 ( .A(n1722), .B(n1377), .Z(n1176) );
  CENX1 U1675 ( .A(n1722), .B(n1376), .Z(n1175) );
  CENX1 U1676 ( .A(n1726), .B(n1377), .Z(n1155) );
  CENX1 U1677 ( .A(n1734), .B(n1378), .Z(n1105) );
  CENX1 U1678 ( .A(n1731), .B(n1376), .Z(n1118) );
  CENX1 U1679 ( .A(n1733), .B(n1377), .Z(n1104) );
  CENX1 U1680 ( .A(n1733), .B(n1376), .Z(n1103) );
  CENX1 U1681 ( .A(n1378), .B(n1738), .Z(n1092) );
  CENX1 U1682 ( .A(n1377), .B(n1738), .Z(n1091) );
  CENX1 U1683 ( .A(n1376), .B(n1738), .Z(n1090) );
  CENX1 U1684 ( .A(n1703), .B(n1378), .Z(n1252) );
  CENX1 U1685 ( .A(n1703), .B(n1377), .Z(n1251) );
  CENX1 U1686 ( .A(n1719), .B(n1378), .Z(n1200) );
  CENX1 U1687 ( .A(n1719), .B(n1376), .Z(n1198) );
  CENX1 U1688 ( .A(n1719), .B(n1377), .Z(n1199) );
  CENX1 U1689 ( .A(n1729), .B(n1377), .Z(n1136) );
  CENX1 U1690 ( .A(n1527), .B(n1378), .Z(n1345) );
  CENX1 U1691 ( .A(n1688), .B(n1377), .Z(n1344) );
  CENX1 U1692 ( .A(n1527), .B(n1376), .Z(n1343) );
  CENX1 U1693 ( .A(n1694), .B(n1371), .Z(n1305) );
  CENX1 U1694 ( .A(n1691), .B(n1378), .Z(n1312) );
  CENX1 U1695 ( .A(n1691), .B(n1377), .Z(n1311) );
  CENX1 U1696 ( .A(n1696), .B(n1377), .Z(n1280) );
  CENX1 U1697 ( .A(n1378), .B(n1740), .Z(n1081) );
  CENX1 U1698 ( .A(n1696), .B(n1378), .Z(n1281) );
  CENX1 U1699 ( .A(n1690), .B(n1376), .Z(n1310) );
  CENX1 U1700 ( .A(n1527), .B(n1375), .Z(n1342) );
  CENX1 U1701 ( .A(n1698), .B(n1376), .Z(n1279) );
  CENX1 U1702 ( .A(n1698), .B(n1375), .Z(n1278) );
  CENX1 U1703 ( .A(n1689), .B(n1371), .Z(n1338) );
  CENX1 U1704 ( .A(n1681), .B(n109), .Z(n1068) );
  CENX1 U1705 ( .A(n104), .B(a[28]), .Z(n110) );
  COND1XL U1706 ( .A(n1674), .B(n1672), .C(n1673), .Z(n286) );
  CENX1 U1707 ( .A(n1726), .B(n1367), .Z(n1145) );
  CENX1 U1708 ( .A(n1719), .B(n1363), .Z(n1185) );
  CENX1 U1709 ( .A(n109), .B(a[30]), .Z(n114) );
  CANR1XL U1710 ( .A(n1678), .B(n286), .C(n283), .Z(n281) );
  CENX1 U1711 ( .A(n1693), .B(b[29]), .Z(n1289) );
  CENX1 U1712 ( .A(n1723), .B(n1365), .Z(n1164) );
  CENX1 U1713 ( .A(n1375), .B(n1738), .Z(n1089) );
  CENX1 U1714 ( .A(n1377), .B(n1740), .Z(n1080) );
  CEOX1 U1715 ( .A(a[4]), .B(n1698), .Z(n1398) );
  CENX1 U1716 ( .A(n1730), .B(n1369), .Z(n1128) );
  CENX1 U1717 ( .A(n1714), .B(n1361), .Z(n1208) );
  CENX1 U1718 ( .A(n1684), .B(n113), .Z(n1066) );
  CENX1 U1719 ( .A(n1686), .B(n113), .Z(n1065) );
  CENX1 U1720 ( .A(n1683), .B(n104), .Z(n1073) );
  CENX1 U1721 ( .A(n1706), .B(n1370), .Z(n1244) );
  CENX1 U1722 ( .A(n1706), .B(n1369), .Z(n1243) );
  CENX1 U1723 ( .A(n1715), .B(n1367), .Z(n1214) );
  CENX1 U1724 ( .A(n1702), .B(n1365), .Z(n1239) );
  CENX1 U1725 ( .A(n1726), .B(n1370), .Z(n1148) );
  CENX1 U1726 ( .A(n1726), .B(n1369), .Z(n1147) );
  CENX1 U1727 ( .A(n1711), .B(n1362), .Z(n1209) );
  CENX1 U1728 ( .A(n1715), .B(n1370), .Z(n1217) );
  CENX1 U1729 ( .A(n1707), .B(n1366), .Z(n1240) );
  CENX1 U1730 ( .A(n1715), .B(n1368), .Z(n1215) );
  CENX1 U1731 ( .A(n1711), .B(n1365), .Z(n1212) );
  CENX1 U1732 ( .A(n1711), .B(n1364), .Z(n1211) );
  CENX1 U1733 ( .A(n1702), .B(n1361), .Z(n1235) );
  CENX1 U1734 ( .A(n1702), .B(n1362), .Z(n1236) );
  CENX1 U1735 ( .A(n1711), .B(n1363), .Z(n1210) );
  CENX1 U1736 ( .A(n1723), .B(n1370), .Z(n1169) );
  CENX1 U1737 ( .A(n1703), .B(n1364), .Z(n1238) );
  CENX1 U1738 ( .A(n1719), .B(n1365), .Z(n1187) );
  CENX1 U1739 ( .A(n1723), .B(n1367), .Z(n1166) );
  CENX1 U1740 ( .A(n1719), .B(n1364), .Z(n1186) );
  CENX1 U1741 ( .A(n1723), .B(n1366), .Z(n1165) );
  CENX1 U1742 ( .A(n1730), .B(n1370), .Z(n1129) );
  CENX1 U1743 ( .A(n1726), .B(n1368), .Z(n1146) );
  CENX1 U1744 ( .A(n1706), .B(n1368), .Z(n1242) );
  CENX1 U1745 ( .A(n1707), .B(n1367), .Z(n1241) );
  CENX1 U1746 ( .A(n1715), .B(n1369), .Z(n1216) );
  CENX1 U1747 ( .A(n1714), .B(n1366), .Z(n1213) );
  CENX1 U1748 ( .A(n1703), .B(n1363), .Z(n1237) );
  CENX1 U1749 ( .A(n1723), .B(n1369), .Z(n1168) );
  CENX1 U1750 ( .A(n1723), .B(n1368), .Z(n1167) );
  CENX1 U1751 ( .A(n1694), .B(n1370), .Z(n1304) );
  CENX1 U1752 ( .A(n1694), .B(n1369), .Z(n1303) );
  CENX1 U1753 ( .A(n1699), .B(n1370), .Z(n1273) );
  CENX1 U1754 ( .A(n1700), .B(n1369), .Z(n1272) );
  CENX1 U1755 ( .A(n1525), .B(n1367), .Z(n1301) );
  CENX1 U1756 ( .A(n1700), .B(n1368), .Z(n1271) );
  CENX1 U1757 ( .A(n1700), .B(n1367), .Z(n1270) );
  CENX1 U1758 ( .A(n1690), .B(n1365), .Z(n1299) );
  CENX1 U1759 ( .A(n1700), .B(n1366), .Z(n1269) );
  CENX1 U1760 ( .A(n1697), .B(n1365), .Z(n1268) );
  CENX1 U1761 ( .A(n1690), .B(n1362), .Z(n1296) );
  CENX1 U1762 ( .A(n1694), .B(n1361), .Z(n1295) );
  CENX1 U1763 ( .A(n1695), .B(n1362), .Z(n1265) );
  CENX1 U1764 ( .A(n1695), .B(n1361), .Z(n1264) );
  CENX1 U1765 ( .A(n1682), .B(n104), .Z(n1074) );
  CENX1 U1766 ( .A(n1690), .B(b[28]), .Z(n1290) );
  CENX1 U1767 ( .A(n1525), .B(n1368), .Z(n1302) );
  CENX1 U1768 ( .A(n1695), .B(n1364), .Z(n1267) );
  CENX1 U1769 ( .A(n1695), .B(n1363), .Z(n1266) );
  CENX1 U1770 ( .A(n1690), .B(b[26]), .Z(n1292) );
  CENX1 U1771 ( .A(n1690), .B(b[27]), .Z(n1291) );
  CENX1 U1772 ( .A(n1689), .B(n1369), .Z(n1336) );
  CENX1 U1773 ( .A(n1689), .B(n1368), .Z(n1335) );
  CENX1 U1774 ( .A(n1688), .B(n1365), .Z(n1332) );
  CENX1 U1775 ( .A(n1690), .B(n1366), .Z(n1300) );
  CENX1 U1776 ( .A(n1688), .B(n1364), .Z(n1331) );
  CENX1 U1777 ( .A(n1688), .B(n1363), .Z(n1330) );
  CENX1 U1778 ( .A(n1691), .B(n1364), .Z(n1298) );
  CENX1 U1779 ( .A(n1691), .B(n1363), .Z(n1297) );
  CENX1 U1780 ( .A(n1688), .B(b[26]), .Z(n1325) );
  CENX1 U1781 ( .A(n1688), .B(b[27]), .Z(n1324) );
  CENX1 U1782 ( .A(n1680), .B(n109), .Z(n1069) );
  CENX1 U1783 ( .A(n1686), .B(n109), .Z(n1070) );
  CENX1 U1784 ( .A(n1688), .B(b[28]), .Z(n1323) );
  CENX1 U1785 ( .A(n1688), .B(b[29]), .Z(n1322) );
  CENX1 U1786 ( .A(n1688), .B(b[30]), .Z(n1321) );
  CENX1 U1787 ( .A(n1689), .B(n1370), .Z(n1337) );
  CENX1 U1788 ( .A(n1689), .B(n1367), .Z(n1334) );
  CENX1 U1789 ( .A(n1527), .B(n1366), .Z(n1333) );
  CENX1 U1790 ( .A(n1688), .B(n1362), .Z(n1329) );
  CENX1 U1791 ( .A(n1688), .B(n1361), .Z(n1328) );
  CENX1 U1792 ( .A(n1681), .B(n104), .Z(n1075) );
  CENX1 U1793 ( .A(n1686), .B(n104), .Z(n1077) );
  CENX1 U1794 ( .A(n1680), .B(n104), .Z(n1076) );
  CENX1 U1795 ( .A(n1527), .B(b[31]), .Z(n1320) );
  CENX1 U1796 ( .A(n1684), .B(n104), .Z(n1078) );
  CENX1 U1797 ( .A(n1684), .B(n109), .Z(n1071) );
  CND2X1 U1798 ( .A(n100), .B(n1388), .Z(n102) );
  CEOXL U1799 ( .A(a[24]), .B(n1740), .Z(n1388) );
  CEOXL U1800 ( .A(a[18]), .B(n1731), .Z(n1391) );
  CNIVX1 U1801 ( .A(n1383), .Z(n1686) );
  CEOXL U1802 ( .A(a[20]), .B(n1734), .Z(n1390) );
  CND2X1 U1803 ( .A(n1387), .B(n105), .Z(n107) );
  CEOXL U1804 ( .A(a[26]), .B(n104), .Z(n1387) );
  CNIVX1 U1805 ( .A(n116), .Z(n1684) );
  CNIVX1 U1806 ( .A(n116), .Z(n1685) );
  COR2X1 U1807 ( .A(n739), .B(n1559), .Z(n1555) );
  CEOXL U1808 ( .A(a[22]), .B(n1738), .Z(n1389) );
  CND2X1 U1809 ( .A(n739), .B(n1559), .Z(n274) );
  CND2X1 U1810 ( .A(n1386), .B(n110), .Z(n112) );
  CEOXL U1811 ( .A(a[28]), .B(n109), .Z(n1386) );
  CEOX1 U1812 ( .A(n1693), .B(a[4]), .Z(n1556) );
  CEOXL U1813 ( .A(a[30]), .B(a[31]), .Z(n1385) );
  CENX1 U1814 ( .A(n142), .B(n286), .Z(product[8]) );
  CND2XL U1815 ( .A(n1678), .B(n1675), .Z(n142) );
  CENX1 U1816 ( .A(n141), .B(n280), .Z(product[9]) );
  CND2XL U1817 ( .A(n334), .B(n1676), .Z(n141) );
  CEOXL U1818 ( .A(n1672), .B(n143), .Z(n1742) );
  CND2XL U1819 ( .A(n336), .B(n1673), .Z(n143) );
  CENX1 U1820 ( .A(n1699), .B(n1371), .Z(n1274) );
  CENX1 U1821 ( .A(n1706), .B(n1371), .Z(n1245) );
  CENX1 U1822 ( .A(n1715), .B(n1371), .Z(n1218) );
  CENX1 U1823 ( .A(n1719), .B(n1371), .Z(n1193) );
  CENX1 U1824 ( .A(n1723), .B(n1371), .Z(n1170) );
  CENX1 U1825 ( .A(n1726), .B(n1371), .Z(n1149) );
  CENX1 U1826 ( .A(n1730), .B(n1371), .Z(n1130) );
  CENX1 U1827 ( .A(n1731), .B(n1371), .Z(n1113) );
  CENX1 U1828 ( .A(n1689), .B(n1372), .Z(n1339) );
  CENX1 U1829 ( .A(n1694), .B(n1372), .Z(n1306) );
  CENX1 U1830 ( .A(n1699), .B(n1372), .Z(n1275) );
  CENX1 U1831 ( .A(n1706), .B(n1372), .Z(n1246) );
  CENX1 U1832 ( .A(n1714), .B(n1372), .Z(n1219) );
  CENX1 U1833 ( .A(n1720), .B(n1372), .Z(n1194) );
  CENX1 U1834 ( .A(n1722), .B(n1372), .Z(n1171) );
  CENX1 U1835 ( .A(n1726), .B(n1372), .Z(n1150) );
  CENX1 U1836 ( .A(n1729), .B(n1372), .Z(n1131) );
  CENXL U1837 ( .A(n1527), .B(n1373), .Z(n1340) );
  CENXL U1838 ( .A(n1693), .B(n1373), .Z(n1307) );
  CENXL U1839 ( .A(n1699), .B(n1373), .Z(n1276) );
  CENXL U1840 ( .A(n1702), .B(n1373), .Z(n1247) );
  CENXL U1841 ( .A(n1715), .B(n1373), .Z(n1220) );
  CENX1 U1842 ( .A(n1726), .B(n1373), .Z(n1151) );
  CENX1 U1843 ( .A(n1730), .B(n1373), .Z(n1132) );
  CENX1 U1844 ( .A(n1731), .B(n1373), .Z(n1115) );
  CENX1 U1845 ( .A(n1734), .B(n1373), .Z(n1100) );
  CENXL U1846 ( .A(n1733), .B(n1375), .Z(n1102) );
  CENXL U1847 ( .A(n1731), .B(n1375), .Z(n1117) );
  CENXL U1848 ( .A(n1729), .B(n1375), .Z(n1134) );
  CENXL U1849 ( .A(n1694), .B(n1375), .Z(n1309) );
  CENXL U1850 ( .A(n1714), .B(n1375), .Z(n1222) );
  CENXL U1851 ( .A(n1722), .B(n1375), .Z(n1174) );
  CENXL U1852 ( .A(n1720), .B(n1375), .Z(n1197) );
  CENXL U1853 ( .A(n1703), .B(n1375), .Z(n1249) );
  CENXL U1854 ( .A(n1726), .B(n1375), .Z(n1153) );
  CENX4 U1855 ( .A(n1527), .B(a[2]), .Z(n15) );
  CND2X4 U1856 ( .A(n1399), .B(n15), .Z(n18) );
  CND2X4 U1857 ( .A(n1398), .B(n24), .Z(n27) );
  CND2X4 U1858 ( .A(n1397), .B(n33), .Z(n36) );
  CND2X4 U1859 ( .A(n1395), .B(n50), .Z(n53) );
  CIVXL U1860 ( .A(n1524), .Z(n1690) );
  CIVXL U1861 ( .A(n1524), .Z(n1691) );
  CIVXL U1862 ( .A(n1524), .Z(n1692) );
  CIVXL U1863 ( .A(n1524), .Z(n1693) );
  CIVXL U1864 ( .A(n1524), .Z(n1694) );
  CIVXL U1865 ( .A(n1701), .Z(n1695) );
  CIVXL U1866 ( .A(n1701), .Z(n1696) );
  CIVXL U1867 ( .A(n1701), .Z(n1697) );
  CIVXL U1868 ( .A(n1701), .Z(n1699) );
  CIVXL U1869 ( .A(n1701), .Z(n1700) );
  CIVXL U1870 ( .A(n1708), .Z(n1702) );
  CIVXL U1871 ( .A(n1709), .Z(n1703) );
  CIVXL U1872 ( .A(n1709), .Z(n1704) );
  CIVXL U1873 ( .A(n1710), .Z(n1706) );
  CIVXL U1874 ( .A(n1710), .Z(n1707) );
  CIVXL U1875 ( .A(n30), .Z(n1708) );
  CIVXL U1876 ( .A(n30), .Z(n1709) );
  CIVXL U1877 ( .A(n30), .Z(n1710) );
  CIVXL U1878 ( .A(n1718), .Z(n1711) );
  CIVXL U1879 ( .A(n1717), .Z(n1712) );
  CIVXL U1880 ( .A(n1717), .Z(n1713) );
  CIVXL U1881 ( .A(n1717), .Z(n1714) );
  CIVXL U1882 ( .A(n1718), .Z(n1715) );
  CIVXL U1883 ( .A(n1718), .Z(n1716) );
  CIVXL U1884 ( .A(n39), .Z(n1717) );
  CIVXL U1885 ( .A(n39), .Z(n1718) );
  CIVX1 U1886 ( .A(n48), .Z(n1721) );
  CIVX1 U1887 ( .A(n55), .Z(n1724) );
  CIVX1 U1888 ( .A(n63), .Z(n1727) );
  CIVXL U1889 ( .A(n79), .Z(n1732) );
  CIVXL U1890 ( .A(n1736), .Z(n1733) );
  CIVXL U1891 ( .A(n1737), .Z(n1734) );
  CIVXL U1892 ( .A(n1737), .Z(n1735) );
  CIVXL U1893 ( .A(n86), .Z(n1736) );
  CIVXL U1894 ( .A(n86), .Z(n1737) );
  CIVX1 U1895 ( .A(n93), .Z(n1739) );
  CIVX1 U1896 ( .A(n99), .Z(n1741) );
  CIVX2 U1897 ( .A(n149), .Z(product[1]) );
  CIVX2 U1898 ( .A(n303), .Z(n340) );
  CIVX2 U1899 ( .A(n295), .Z(n338) );
  CIVX2 U1900 ( .A(n1674), .Z(n336) );
  CIVX2 U1901 ( .A(n265), .Z(n332) );
  CIVX2 U1902 ( .A(n262), .Z(n331) );
  CIVX2 U1903 ( .A(n224), .Z(n325) );
  CIVX2 U1904 ( .A(n159), .Z(n315) );
  CIVX2 U1905 ( .A(n151), .Z(n313) );
  CIVX2 U1906 ( .A(n312), .Z(n310) );
  CIVX2 U1907 ( .A(n309), .Z(n307) );
  CIVX2 U1908 ( .A(n301), .Z(n299) );
  CIVX2 U1909 ( .A(n293), .Z(n291) );
  CIVX2 U1910 ( .A(n1675), .Z(n283) );
  CIVX2 U1911 ( .A(n281), .Z(n280) );
  CIVX2 U1912 ( .A(n1676), .Z(n277) );
  CIVX2 U1913 ( .A(n1677), .Z(n334) );
  CIVX2 U1914 ( .A(n274), .Z(n272) );
  CIVX2 U1915 ( .A(n268), .Z(n267) );
  CIVX2 U1916 ( .A(n259), .Z(n258) );
  CIVX2 U1917 ( .A(n257), .Z(n255) );
  CIVX2 U1918 ( .A(n256), .Z(n330) );
  CIVX2 U1919 ( .A(n247), .Z(n245) );
  CIVX2 U1920 ( .A(n235), .Z(n237) );
  CIVX2 U1921 ( .A(n234), .Z(n327) );
  CIVX2 U1922 ( .A(n232), .Z(n230) );
  CIVX2 U1923 ( .A(n219), .Z(n217) );
  CIVX2 U1924 ( .A(n214), .Z(n212) );
  CIVX2 U1925 ( .A(n192), .Z(n190) );
  CIVX2 U1926 ( .A(n187), .Z(n185) );
  CIVX2 U1927 ( .A(n177), .Z(n175) );
  CIVX2 U1928 ( .A(n172), .Z(n170) );
  CIVX2 U1929 ( .A(n165), .Z(n163) );
  CIVX2 U1930 ( .A(n157), .Z(n155) );
  CIVX2 U1931 ( .A(n104), .Z(n1412) );
  CIVX2 U1932 ( .A(n109), .Z(n1411) );
  CIVX2 U1933 ( .A(n113), .Z(n1410) );
endmodule


module calc_DW02_mult_2_stage_7 ( A, B, TC, CLK, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC, CLK;
  wire   n26, n27, n28, n29, n30, n31, n32, \A_extended[32] , \B_extended[32] ,
         n6, n8, n10, n12, n14, n16, n18, n19, n20, n21, n22, n23, n24, n25;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33;
  assign \A_extended[32]  = A[31];
  assign \B_extended[32]  = B[31];

  calc_DW_mult_tc_17 mult_96 ( .a({\A_extended[32] , \A_extended[32] , A[30:0]}), .b({\B_extended[32] , \B_extended[32] , B[30:0]}), .product({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, PRODUCT[31:7], n26, 
        n27, n28, n29, n30, n31, n32}), .dw4_CLK(CLK) );
  CFD1QXL clk_r_REG127_S1 ( .D(n32), .CP(CLK), .Q(n19) );
  CFD1QXL clk_r_REG126_S1 ( .D(n31), .CP(CLK), .Q(n20) );
  CFD1QXL clk_r_REG119_S1 ( .D(n26), .CP(CLK), .Q(n25) );
  CFD1QXL clk_r_REG121_S1 ( .D(n27), .CP(CLK), .Q(n24) );
  CFD1QXL clk_r_REG123_S1 ( .D(n28), .CP(CLK), .Q(n23) );
  CFD1QXL clk_r_REG124_S1 ( .D(n29), .CP(CLK), .Q(n22) );
  CFD1QXL clk_r_REG125_S1 ( .D(n30), .CP(CLK), .Q(n21) );
  CIVDXL U1 ( .A(n24), .Z1(n6) );
  CNIVX1 U2 ( .A(n6), .Z(PRODUCT[5]) );
  CIVDXL U3 ( .A(n19), .Z1(n8) );
  CNIVX1 U4 ( .A(n8), .Z(PRODUCT[0]) );
  CIVDXL U5 ( .A(n22), .Z1(n10) );
  CNIVX1 U6 ( .A(n10), .Z(PRODUCT[3]) );
  CIVDXL U7 ( .A(n21), .Z1(n12) );
  CNIVX1 U8 ( .A(n12), .Z(PRODUCT[2]) );
  CIVDXL U9 ( .A(n20), .Z1(n14) );
  CNIVX1 U10 ( .A(n14), .Z(PRODUCT[1]) );
  CIVDXL U11 ( .A(n25), .Z1(n16) );
  CNIVX1 U12 ( .A(n16), .Z(PRODUCT[6]) );
  CIVDXL U13 ( .A(n23), .Z1(n18) );
  CNIVX1 U14 ( .A(n18), .Z(PRODUCT[4]) );
endmodule


module calc_DW_mult_tc_19 ( a, b, product, dw3_CLK );
  input [32:0] a;
  input [32:0] b;
  output [65:0] product;
  input dw3_CLK;
  wire   n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n32, n34, n36, n38, n40, n42, n44, n46, n48, n50, n52, n54,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n90, n92, n93, n94, n95, n96, n98, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n117,
         n118, n119, n120, n122, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n135, n137, n138, n139, n140, n142, n145, n146,
         n147, n148, n150, n152, n153, n155, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n172, n174,
         n175, n177, n179, n180, n181, n183, n185, n186, n187, n188, n189,
         n191, n193, n194, n195, n196, n197, n199, n201, n202, n203, n204,
         n205, n207, n209, n210, n212, n213, n216, n218, n219, n220, n221,
         n223, n225, n229, n233, n235, n237, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n885, n910, n911, n912, \b[0] , n1094, n1093, n1092, n1091,
         n986, n988, n990, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060;
  assign product[0] = \b[0] ;
  assign \b[0]  = b[0];
  assign n1060 = dw3_CLK;

  CFA1X1 U50 ( .A(n282), .B(n86), .CI(n255), .CO(n85), .S(product[30]) );
  CFA1X1 U51 ( .A(n308), .B(n87), .CI(n283), .CO(n86), .S(product[29]) );
  CFA1X1 U52 ( .A(n334), .B(n1005), .CI(n309), .CO(n87), .S(product[28]) );
  CEO3X2 U257 ( .A(n260), .B(n243), .C(n242), .Z(n241) );
  CEO3X2 U258 ( .A(n245), .B(n262), .C(n244), .Z(n242) );
  CEO3X2 U259 ( .A(n246), .B(n247), .C(n264), .Z(n243) );
  CEO3X2 U260 ( .A(n248), .B(n268), .C(n266), .Z(n244) );
  CEO3X2 U261 ( .A(n249), .B(n250), .C(n270), .Z(n245) );
  CEO3X2 U262 ( .A(n274), .B(n251), .C(n252), .Z(n246) );
  CEO3X2 U263 ( .A(n276), .B(n272), .C(n253), .Z(n247) );
  CEO3X2 U266 ( .A(n667), .B(n674), .C(n682), .Z(n250) );
  CEO3X2 U268 ( .A(n701), .B(n649), .C(n751), .Z(n252) );
  CFA1X1 U270 ( .A(n1028), .B(n1029), .CI(n1027), .CO(n254), .S(n255) );
  CFA1X1 U271 ( .A(n288), .B(n286), .CI(n261), .CO(n256), .S(n257) );
  CFA1X1 U272 ( .A(n265), .B(n263), .CI(n290), .CO(n258), .S(n259) );
  CFA1X1 U273 ( .A(n269), .B(n267), .CI(n292), .CO(n260), .S(n261) );
  CFA1X1 U274 ( .A(n271), .B(n294), .CI(n296), .CO(n262), .S(n263) );
  CFA1X1 U275 ( .A(n275), .B(n277), .CI(n273), .CO(n264), .S(n265) );
  CFA1X1 U276 ( .A(n298), .B(n279), .CI(n300), .CO(n266), .S(n267) );
  CFA1X1 U277 ( .A(n281), .B(n302), .CI(n304), .CO(n268), .S(n269) );
  CFA1X1 U278 ( .A(n692), .B(n306), .CI(n713), .CO(n270), .S(n271) );
  CFA1X1 U279 ( .A(n725), .B(n683), .CI(n657), .CO(n272), .S(n273) );
  CFA1X1 U281 ( .A(n675), .B(n752), .CI(n650), .CO(n276), .S(n277) );
  CFA1X1 U282 ( .A(n702), .B(n766), .CI(n648), .CO(n278), .S(n279) );
  CHA1X1 U283 ( .A(a[15]), .B(n662), .CO(n280), .S(n281) );
  CFA1X1 U284 ( .A(n1025), .B(n1026), .CI(n1024), .CO(n282), .S(n283) );
  CFA1X1 U285 ( .A(n291), .B(n312), .CI(n289), .CO(n284), .S(n285) );
  CFA1X1 U286 ( .A(n316), .B(n314), .CI(n293), .CO(n286), .S(n287) );
  CFA1X1 U287 ( .A(n297), .B(n295), .CI(n318), .CO(n288), .S(n289) );
  CFA1X1 U288 ( .A(n301), .B(n320), .CI(n299), .CO(n290), .S(n291) );
  CFA1X1 U289 ( .A(n305), .B(n322), .CI(n303), .CO(n292), .S(n293) );
  CFA1X1 U290 ( .A(n328), .B(n326), .CI(n324), .CO(n294), .S(n295) );
  CFA1X1 U291 ( .A(n332), .B(n330), .CI(n307), .CO(n296), .S(n297) );
  CFA1X1 U292 ( .A(n714), .B(n693), .CI(n676), .CO(n298), .S(n299) );
  CFA1X1 U294 ( .A(n684), .B(n739), .CI(n753), .CO(n302), .S(n303) );
  CFA1X1 U295 ( .A(n703), .B(n654), .CI(n767), .CO(n304), .S(n305) );
  CHA1X1 U296 ( .A(n663), .B(n651), .CO(n306), .S(n307) );
  CFA1X1 U297 ( .A(n1022), .B(n1023), .CI(n1021), .CO(n308), .S(n309) );
  CFA1X1 U298 ( .A(n340), .B(n338), .CI(n315), .CO(n310), .S(n311) );
  CFA1X1 U299 ( .A(n342), .B(n317), .CI(n319), .CO(n312), .S(n313) );
  CFA1X1 U300 ( .A(n346), .B(n321), .CI(n344), .CO(n314), .S(n315) );
  CFA1X1 U301 ( .A(n331), .B(n323), .CI(n329), .CO(n316), .S(n317) );
  CFA1X1 U302 ( .A(n348), .B(n325), .CI(n327), .CO(n318), .S(n319) );
  CFA1X1 U303 ( .A(n354), .B(n352), .CI(n350), .CO(n320), .S(n321) );
  CFA1X1 U304 ( .A(n715), .B(n333), .CI(n356), .CO(n322), .S(n323) );
  CFA1X1 U305 ( .A(n727), .B(n694), .CI(n677), .CO(n324), .S(n325) );
  CFA1X1 U306 ( .A(n670), .B(n659), .CI(n740), .CO(n326), .S(n327) );
  CFA1X1 U307 ( .A(n685), .B(n754), .CI(n655), .CO(n328), .S(n329) );
  CFA1X1 U308 ( .A(n664), .B(n781), .CI(n768), .CO(n330), .S(n331) );
  CHA1X1 U309 ( .A(a[14]), .B(n704), .CO(n332), .S(n333) );
  CFA1X1 U310 ( .A(n1019), .B(n1020), .CI(n1018), .CO(n334), .S(n335) );
  CFA1X1 U311 ( .A(n364), .B(n362), .CI(n341), .CO(n336), .S(n337) );
  CFA1X1 U312 ( .A(n366), .B(n343), .CI(n345), .CO(n338), .S(n339) );
  CFA1X1 U313 ( .A(n370), .B(n347), .CI(n368), .CO(n340), .S(n341) );
  CFA1X1 U314 ( .A(n353), .B(n349), .CI(n351), .CO(n342), .S(n343) );
  CFA1X1 U315 ( .A(n374), .B(n355), .CI(n372), .CO(n344), .S(n345) );
  CFA1X1 U316 ( .A(n357), .B(n376), .CI(n378), .CO(n346), .S(n347) );
  CFA1X1 U317 ( .A(n741), .B(n380), .CI(n728), .CO(n348), .S(n349) );
  CFA1X1 U318 ( .A(n755), .B(n716), .CI(n695), .CO(n350), .S(n351) );
  CFA1X1 U320 ( .A(n705), .B(n660), .CI(n769), .CO(n354), .S(n355) );
  CHA1X1 U321 ( .A(n665), .B(n782), .CO(n356), .S(n357) );
  CFA1X1 U322 ( .A(n1016), .B(n1017), .CI(n1013), .CO(n358), .S(n359) );
  CFA1X1 U323 ( .A(n388), .B(n386), .CI(n365), .CO(n360), .S(n361) );
  CFA1X1 U324 ( .A(n390), .B(n367), .CI(n369), .CO(n362), .S(n363) );
  CFA1X1 U325 ( .A(n394), .B(n371), .CI(n392), .CO(n364), .S(n365) );
  CFA1X1 U326 ( .A(n373), .B(n375), .CI(n377), .CO(n366), .S(n367) );
  CFA1X1 U327 ( .A(n398), .B(n379), .CI(n396), .CO(n368), .S(n369) );
  CFA1X1 U328 ( .A(n402), .B(n400), .CI(n381), .CO(n370), .S(n371) );
  CFA1X1 U329 ( .A(n756), .B(n742), .CI(n729), .CO(n372), .S(n373) );
  CFA1X1 U330 ( .A(n770), .B(n717), .CI(n687), .CO(n374), .S(n375) );
  CFA1X1 U331 ( .A(n696), .B(n679), .CI(n672), .CO(n376), .S(n377) );
  CFA1X1 U332 ( .A(n706), .B(n783), .CI(n795), .CO(n378), .S(n379) );
  CHA1X1 U333 ( .A(a[13]), .B(n666), .CO(n380), .S(n381) );
  CFA1X1 U334 ( .A(n387), .B(n385), .CI(n406), .CO(n382), .S(n383) );
  CFA1X1 U335 ( .A(n391), .B(n389), .CI(n408), .CO(n384), .S(n385) );
  CFA1X1 U336 ( .A(n412), .B(n410), .CI(n393), .CO(n386), .S(n387) );
  CFA1X1 U337 ( .A(n397), .B(n395), .CI(n414), .CO(n388), .S(n389) );
  CFA1X1 U338 ( .A(n416), .B(n399), .CI(n401), .CO(n390), .S(n391) );
  CFA1X1 U339 ( .A(n422), .B(n420), .CI(n418), .CO(n392), .S(n393) );
  CFA1X1 U340 ( .A(n743), .B(n403), .CI(n424), .CO(n394), .S(n395) );
  CFA1X1 U341 ( .A(n757), .B(n697), .CI(n688), .CO(n396), .S(n397) );
  CFA1X1 U342 ( .A(n730), .B(n771), .CI(n784), .CO(n398), .S(n399) );
  CFA1X1 U343 ( .A(n718), .B(n680), .CI(n673), .CO(n400), .S(n401) );
  CHA1X1 U344 ( .A(n707), .B(n796), .CO(n402), .S(n403) );
  CFA1X1 U345 ( .A(n409), .B(n407), .CI(n428), .CO(n404), .S(n405) );
  CFA1X1 U346 ( .A(n413), .B(n430), .CI(n411), .CO(n406), .S(n407) );
  CFA1X1 U347 ( .A(n434), .B(n432), .CI(n415), .CO(n408), .S(n409) );
  CFA1X1 U348 ( .A(n423), .B(n436), .CI(n417), .CO(n410), .S(n411) );
  CFA1X1 U349 ( .A(n438), .B(n421), .CI(n419), .CO(n412), .S(n413) );
  CFA1X1 U350 ( .A(n425), .B(n440), .CI(n442), .CO(n414), .S(n415) );
  CFA1X1 U351 ( .A(n731), .B(n444), .CI(n719), .CO(n416), .S(n417) );
  CFA1X1 U352 ( .A(n758), .B(n689), .CI(n681), .CO(n418), .S(n419) );
  CFA1X1 U353 ( .A(n698), .B(n772), .CI(n797), .CO(n420), .S(n421) );
  CFA1X1 U354 ( .A(n744), .B(n785), .CI(n808), .CO(n422), .S(n423) );
  CHA1X1 U355 ( .A(a[12]), .B(n708), .CO(n424), .S(n425) );
  CFA1X1 U356 ( .A(n431), .B(n429), .CI(n448), .CO(n426), .S(n427) );
  CFA1X1 U357 ( .A(n435), .B(n450), .CI(n433), .CO(n428), .S(n429) );
  CFA1X1 U358 ( .A(n454), .B(n452), .CI(n437), .CO(n430), .S(n431) );
  CFA1X1 U359 ( .A(n443), .B(n456), .CI(n441), .CO(n432), .S(n433) );
  CFA1X1 U360 ( .A(n460), .B(n439), .CI(n458), .CO(n434), .S(n435) );
  CFA1X1 U361 ( .A(n464), .B(n462), .CI(n445), .CO(n436), .S(n437) );
  CFA1X1 U362 ( .A(n773), .B(n759), .CI(n745), .CO(n438), .S(n439) );
  CFA1X1 U363 ( .A(n720), .B(n699), .CI(n690), .CO(n440), .S(n441) );
  CFA1X1 U364 ( .A(n732), .B(n786), .CI(n809), .CO(n442), .S(n443) );
  CHA1X1 U365 ( .A(n709), .B(n798), .CO(n444), .S(n445) );
  CFA1X1 U366 ( .A(n451), .B(n449), .CI(n468), .CO(n446), .S(n447) );
  CFA1X1 U367 ( .A(n455), .B(n470), .CI(n453), .CO(n448), .S(n449) );
  CFA1X1 U368 ( .A(n457), .B(n472), .CI(n474), .CO(n450), .S(n451) );
  CFA1X1 U369 ( .A(n459), .B(n461), .CI(n463), .CO(n452), .S(n453) );
  CFA1X1 U370 ( .A(n480), .B(n476), .CI(n478), .CO(n454), .S(n455) );
  CFA1X1 U371 ( .A(n746), .B(n465), .CI(n482), .CO(n456), .S(n457) );
  CFA1X1 U372 ( .A(n760), .B(n721), .CI(n700), .CO(n458), .S(n459) );
  CFA1X1 U373 ( .A(n733), .B(n787), .CI(n774), .CO(n460), .S(n461) );
  CFA1X1 U374 ( .A(n820), .B(n799), .CI(n810), .CO(n462), .S(n463) );
  CHA1X1 U375 ( .A(a[11]), .B(n710), .CO(n464), .S(n465) );
  CFA1X1 U376 ( .A(n471), .B(n469), .CI(n486), .CO(n466), .S(n467) );
  CFA1X1 U377 ( .A(n490), .B(n488), .CI(n473), .CO(n468), .S(n469) );
  CFA1X1 U378 ( .A(n477), .B(n475), .CI(n492), .CO(n470), .S(n471) );
  CFA1X1 U379 ( .A(n494), .B(n481), .CI(n479), .CO(n472), .S(n473) );
  CFA1X1 U380 ( .A(n483), .B(n496), .CI(n498), .CO(n474), .S(n475) );
  CFA1X1 U381 ( .A(n775), .B(n500), .CI(n747), .CO(n476), .S(n477) );
  CFA1X1 U382 ( .A(n734), .B(n811), .CI(n722), .CO(n478), .S(n479) );
  CFA1X1 U383 ( .A(n761), .B(n800), .CI(n788), .CO(n480), .S(n481) );
  CHA1X1 U384 ( .A(n711), .B(n821), .CO(n482), .S(n483) );
  CFA1X1 U385 ( .A(n489), .B(n487), .CI(n504), .CO(n484), .S(n485) );
  CFA1X1 U386 ( .A(n493), .B(n506), .CI(n491), .CO(n486), .S(n487) );
  CFA1X1 U387 ( .A(n499), .B(n508), .CI(n510), .CO(n488), .S(n489) );
  CFA1X1 U388 ( .A(n512), .B(n497), .CI(n495), .CO(n490), .S(n491) );
  CFA1X1 U389 ( .A(n516), .B(n514), .CI(n501), .CO(n492), .S(n493) );
  CFA1X1 U390 ( .A(n789), .B(n776), .CI(n748), .CO(n494), .S(n495) );
  CFA1X1 U391 ( .A(n762), .B(n822), .CI(n723), .CO(n496), .S(n497) );
  CFA1X1 U392 ( .A(n831), .B(n801), .CI(n812), .CO(n498), .S(n499) );
  CHA1X1 U393 ( .A(a[10]), .B(n735), .CO(n500), .S(n501) );
  CFA1X1 U394 ( .A(n507), .B(n505), .CI(n520), .CO(n502), .S(n503) );
  CFA1X1 U395 ( .A(n511), .B(n509), .CI(n522), .CO(n504), .S(n505) );
  CFA1X1 U396 ( .A(n513), .B(n524), .CI(n515), .CO(n506), .S(n507) );
  CFA1X1 U397 ( .A(n530), .B(n526), .CI(n528), .CO(n508), .S(n509) );
  CFA1X1 U398 ( .A(n832), .B(n517), .CI(n532), .CO(n510), .S(n511) );
  CFA1X1 U399 ( .A(n986), .B(n802), .CI(n994), .CO(n512), .S(n513) );
  CFA1X1 U400 ( .A(n777), .B(n823), .CI(n813), .CO(n514), .S(n515) );
  CHA1X1 U401 ( .A(n736), .B(n790), .CO(n516), .S(n517) );
  CFA1X1 U402 ( .A(n523), .B(n521), .CI(n536), .CO(n518), .S(n519) );
  CFA1X1 U403 ( .A(n540), .B(n538), .CI(n525), .CO(n520), .S(n521) );
  CFA1X1 U404 ( .A(n529), .B(n527), .CI(n531), .CO(n522), .S(n523) );
  CFA1X1 U405 ( .A(n533), .B(n542), .CI(n544), .CO(n524), .S(n525) );
  CFA1X1 U406 ( .A(n833), .B(n546), .CI(n764), .CO(n526), .S(n527) );
  CFA1X1 U407 ( .A(n778), .B(n791), .CI(n824), .CO(n528), .S(n529) );
  CFA1X1 U408 ( .A(n814), .B(n841), .CI(n803), .CO(n530), .S(n531) );
  CHA1X1 U409 ( .A(a[9]), .B(n750), .CO(n532), .S(n533) );
  CFA1X1 U410 ( .A(n539), .B(n537), .CI(n550), .CO(n534), .S(n535) );
  CFA1X1 U411 ( .A(n554), .B(n552), .CI(n541), .CO(n536), .S(n537) );
  CFA1X1 U412 ( .A(n556), .B(n545), .CI(n543), .CO(n538), .S(n539) );
  CFA1X1 U413 ( .A(n560), .B(n558), .CI(n547), .CO(n540), .S(n541) );
  CFA1X1 U414 ( .A(n825), .B(n804), .CI(n765), .CO(n542), .S(n543) );
  CFA1X1 U415 ( .A(n834), .B(n792), .CI(n842), .CO(n544), .S(n545) );
  CHA1X1 U416 ( .A(n779), .B(n815), .CO(n546), .S(n547) );
  CFA1X1 U417 ( .A(n553), .B(n551), .CI(n564), .CO(n548), .S(n549) );
  CFA1X1 U418 ( .A(n557), .B(n566), .CI(n555), .CO(n550), .S(n551) );
  CFA1X1 U419 ( .A(n570), .B(n559), .CI(n568), .CO(n552), .S(n553) );
  CFA1X1 U420 ( .A(n843), .B(n561), .CI(n572), .CO(n554), .S(n555) );
  CFA1X1 U421 ( .A(n816), .B(n826), .CI(n850), .CO(n556), .S(n557) );
  CFA1X1 U422 ( .A(n835), .B(n805), .CI(n793), .CO(n558), .S(n559) );
  CHA1X1 U423 ( .A(a[8]), .B(n780), .CO(n560), .S(n561) );
  CFA1X1 U424 ( .A(n567), .B(n565), .CI(n576), .CO(n562), .S(n563) );
  CFA1X1 U425 ( .A(n571), .B(n578), .CI(n569), .CO(n564), .S(n565) );
  CFA1X1 U426 ( .A(n573), .B(n580), .CI(n582), .CO(n566), .S(n567) );
  CFA1X1 U427 ( .A(n817), .B(n584), .CI(n806), .CO(n568), .S(n569) );
  CFA1X1 U428 ( .A(n836), .B(n827), .CI(n851), .CO(n570), .S(n571) );
  CHA1X1 U429 ( .A(n844), .B(n794), .CO(n572), .S(n573) );
  CFA1X1 U430 ( .A(n579), .B(n577), .CI(n588), .CO(n574), .S(n575) );
  CFA1X1 U431 ( .A(n583), .B(n590), .CI(n581), .CO(n576), .S(n577) );
  CFA1X1 U432 ( .A(n594), .B(n592), .CI(n585), .CO(n578), .S(n579) );
  CFA1X1 U433 ( .A(n845), .B(n828), .CI(n818), .CO(n580), .S(n581) );
  CFA1X1 U434 ( .A(n837), .B(n858), .CI(n807), .CO(n582), .S(n583) );
  CHA1X1 U435 ( .A(a[7]), .B(n852), .CO(n584), .S(n585) );
  CFA1X1 U436 ( .A(n591), .B(n589), .CI(n598), .CO(n586), .S(n587) );
  CFA1X1 U437 ( .A(n602), .B(n593), .CI(n600), .CO(n588), .S(n589) );
  CFA1X1 U438 ( .A(n846), .B(n595), .CI(n604), .CO(n590), .S(n591) );
  CFA1X1 U439 ( .A(n859), .B(n829), .CI(n853), .CO(n592), .S(n593) );
  CHA1X1 U440 ( .A(n838), .B(n819), .CO(n594), .S(n595) );
  CFA1X1 U441 ( .A(n601), .B(n599), .CI(n608), .CO(n596), .S(n597) );
  CFA1X1 U442 ( .A(n605), .B(n603), .CI(n610), .CO(n598), .S(n599) );
  CFA1X1 U443 ( .A(n854), .B(n612), .CI(n847), .CO(n600), .S(n601) );
  CFA1X1 U444 ( .A(n865), .B(n860), .CI(n830), .CO(n602), .S(n603) );
  CHA1X1 U445 ( .A(a[6]), .B(n839), .CO(n604), .S(n605) );
  CFA1X1 U446 ( .A(n611), .B(n609), .CI(n616), .CO(n606), .S(n607) );
  CFA1X1 U447 ( .A(n620), .B(n618), .CI(n613), .CO(n608), .S(n609) );
  CFA1X1 U448 ( .A(n855), .B(n866), .CI(n861), .CO(n610), .S(n611) );
  CHA1X1 U449 ( .A(n840), .B(n848), .CO(n612), .S(n613) );
  CFA1X1 U450 ( .A(n624), .B(n617), .CI(n619), .CO(n614), .S(n615) );
  CFA1X1 U451 ( .A(n862), .B(n621), .CI(n626), .CO(n616), .S(n617) );
  CFA1X1 U452 ( .A(n867), .B(n856), .CI(n849), .CO(n618), .S(n619) );
  CHA1X1 U453 ( .A(a[5]), .B(n871), .CO(n620), .S(n621) );
  CFA1X1 U454 ( .A(n627), .B(n625), .CI(n630), .CO(n622), .S(n623) );
  CFA1X1 U455 ( .A(n868), .B(n632), .CI(n863), .CO(n624), .S(n625) );
  CHA1X1 U456 ( .A(n872), .B(n857), .CO(n626), .S(n627) );
  CFA1X1 U457 ( .A(n636), .B(n631), .CI(n633), .CO(n628), .S(n629) );
  CFA1X1 U458 ( .A(n876), .B(n869), .CI(n864), .CO(n630), .S(n631) );
  CHA1X1 U459 ( .A(a[4]), .B(n873), .CO(n632), .S(n633) );
  CFA1X1 U460 ( .A(n877), .B(n637), .CI(n640), .CO(n634), .S(n635) );
  CHA1X1 U461 ( .A(n874), .B(n870), .CO(n636), .S(n637) );
  CFA1X1 U462 ( .A(n880), .B(n642), .CI(n878), .CO(n638), .S(n639) );
  CHA1X1 U463 ( .A(a[3]), .B(n875), .CO(n640), .S(n641) );
  CHA1X1 U464 ( .A(n881), .B(n879), .CO(n642), .S(n643) );
  CFD1QXL clk_r_REG49_S1 ( .D(n998), .CP(n1060), .Q(n1055) );
  CFD1QXL clk_r_REG48_S1 ( .D(n177), .CP(n1060), .Q(n1054) );
  CFD1QXL clk_r_REG0_S1 ( .D(n257), .CP(n1060), .Q(n1029) );
  CFD1QXL clk_r_REG44_S1 ( .D(n165), .CP(n1060), .Q(n1036) );
  CFD1QXL clk_r_REG43_S1 ( .D(n166), .CP(n1060), .Q(n1035) );
  CFD1QXL clk_r_REG3_S1 ( .D(n284), .CP(n1060), .Q(n1027) );
  CFD1QXL clk_r_REG6_S1 ( .D(n259), .CP(n1060), .Q(n1028) );
  CFD1QXL clk_r_REG36_S1 ( .D(n73), .CP(n1060), .Q(n1037) );
  CFD1QXL clk_r_REG41_S1 ( .D(n75), .CP(n1060), .Q(n1034) );
  CFD1QXL clk_r_REG47_S1 ( .D(n76), .CP(n1060), .Q(n1033) );
  CFD1QXL clk_r_REG1_S1 ( .D(n240), .CP(n1060), .Q(n1030) );
  CFD1QXL clk_r_REG46_S1 ( .D(n180), .CP(n1060), .Q(n1053) );
  CFD1QXL clk_r_REG38_S1 ( .D(n160), .CP(n1060), .Q(n1038) );
  CFD1QXL clk_r_REG37_S1 ( .D(n161), .CP(n1060), .Q(n1032) );
  CFD1QXL clk_r_REG4_S1 ( .D(n285), .CP(n1060), .Q(n1026) );
  CFD1QXL clk_r_REG42_S1 ( .D(n168), .CP(n1060), .Q(n1031) );
  CFD1QXL clk_r_REG35_S1 ( .D(n139), .CP(n1060), .Q(n1042) );
  CFD1QXL clk_r_REG21_S1 ( .D(n108), .CP(n1060), .Q(n1051) );
  CFD1QXL clk_r_REG11_S1 ( .D(n310), .CP(n1060), .Q(n1024) );
  CFD1QXL clk_r_REG9_S1 ( .D(n336), .CP(n1060), .Q(n1021) );
  CFD1QXL clk_r_REG7_S1 ( .D(n360), .CP(n1060), .Q(n1018) );
  CFD1QXL clk_r_REG16_S1 ( .D(n384), .CP(n1060), .Q(n1013) );
  CFD1QXL clk_r_REG5_S1 ( .D(n287), .CP(n1060), .Q(n1025) );
  CFD1QXL clk_r_REG2_S1 ( .D(n313), .CP(n1060), .Q(n1022) );
  CFD1QXL clk_r_REG13_S1 ( .D(n339), .CP(n1060), .Q(n1019) );
  CFD1QXL clk_r_REG58_S1 ( .D(n363), .CP(n1060), .Q(n1016) );
  CFD1QXL clk_r_REG32_S1 ( .D(n152), .CP(n1060), .Q(n1040) );
  CFD1QXL clk_r_REG28_S1 ( .D(n137), .CP(n1060), .Q(n1043) );
  CFD1QXL clk_r_REG39_S1 ( .D(n157), .CP(n1060), .Q(n1039) );
  CFD1QXL clk_r_REG18_S1 ( .D(n383), .CP(n1060), .Q(n1014) );
  CFD1QXL clk_r_REG15_S1 ( .D(n405), .CP(n1060), .Q(n1011) );
  CFD1QXL clk_r_REG19_S1 ( .D(n111), .CP(n1060), .Q(n1049) );
  CFD1QXL clk_r_REG17_S1 ( .D(n382), .CP(n1060), .Q(n1015) );
  CFD1QXL clk_r_REG14_S1 ( .D(n404), .CP(n1060), .Q(n1012) );
  CFD1QXL clk_r_REG23_S1 ( .D(n426), .CP(n1060), .Q(n1010) );
  CFD1QXL clk_r_REG22_S1 ( .D(n107), .CP(n1060), .Q(n1052) );
  CFD1QXL clk_r_REG33_S1 ( .D(n995), .CP(n1060), .Q(n1057) );
  CFD1QXL clk_r_REG29_S1 ( .D(n996), .CP(n1060), .Q(n1058) );
  CFD1QXL clk_r_REG20_S1 ( .D(n110), .CP(n1060), .Q(n1050) );
  CFD1QXL clk_r_REG34_S1 ( .D(n140), .CP(n1060), .Q(n1041) );
  CFD1QXL clk_r_REG25_S1 ( .D(n997), .CP(n1060), .Q(n1059) );
  CFD1QXL clk_r_REG40_S1 ( .D(n1001), .CP(n1060), .Q(n1056) );
  CFD1QXL clk_r_REG8_S1 ( .D(n361), .CP(n1060), .Q(n1017) );
  CFD1QXL clk_r_REG12_S1 ( .D(n311), .CP(n1060), .Q(n1023) );
  CFD1QXL clk_r_REG27_S1 ( .D(n118), .CP(n1060), .Q(n1048) );
  CFD1QXL clk_r_REG24_S1 ( .D(n124), .CP(n1060), .Q(n1046) );
  CFD1QXL clk_r_REG30_S1 ( .D(n130), .CP(n1060), .Q(n1044) );
  CFD1QXL clk_r_REG31_S1 ( .D(n129), .CP(n1060), .Q(n1045) );
  CFD1QXL clk_r_REG26_S1 ( .D(n119), .CP(n1060), .Q(n1047) );
  CFD1QXL clk_r_REG10_S1 ( .D(n337), .CP(n1060), .Q(n1020) );
  CEO3X1 U754 ( .A(n258), .B(n241), .C(n256), .Z(n240) );
  CIVXL U755 ( .A(n113), .Z(n112) );
  CANR1X2 U756 ( .A(n1009), .B(n101), .C(n98), .Z(n96) );
  CIVX2 U757 ( .A(b[17]), .Z(n17) );
  COND1X1 U758 ( .A(n94), .B(n96), .C(n95), .Z(n93) );
  CNIVX1 U759 ( .A(n749), .Z(n986) );
  CIVX8 U760 ( .A(\b[0] ), .Z(n32) );
  CNR2X1 U761 ( .A(n32), .B(n20), .Z(n711) );
  CNR2X1 U762 ( .A(n32), .B(n17), .Z(n750) );
  CND2XL U763 ( .A(n220), .B(n1049), .Z(n65) );
  CIVXL U764 ( .A(n159), .Z(n158) );
  CNIVX1 U765 ( .A(n988), .Z(product[11]) );
  CNIVX1 U766 ( .A(n1094), .Z(n988) );
  CNIVX1 U767 ( .A(n990), .Z(product[12]) );
  CNIVX1 U768 ( .A(n1093), .Z(n990) );
  CNIVX1 U769 ( .A(n1092), .Z(product[13]) );
  CNIVX1 U770 ( .A(n993), .Z(product[14]) );
  CNIVX1 U771 ( .A(n1091), .Z(n993) );
  CFA1XL U772 ( .A(n668), .B(n653), .CI(n738), .CO(n274), .S(n275) );
  CANR1X1 U773 ( .A(n1038), .B(n1031), .C(n1032), .Z(n159) );
  COND1X1 U774 ( .A(n147), .B(n159), .C(n148), .Z(n146) );
  CANR1X1 U775 ( .A(n155), .B(n1057), .C(n150), .Z(n148) );
  CENXL U776 ( .A(n93), .B(n60), .Z(product[27]) );
  CHA1XL U777 ( .A(a[2]), .B(n883), .CO(n644), .S(n645) );
  CIVX4 U778 ( .A(b[2]), .Z(n36) );
  CFA1XL U779 ( .A(n726), .B(n669), .CI(n658), .CO(n300), .S(n301) );
  CNR2X1 U780 ( .A(n36), .B(n26), .Z(n658) );
  CFA1XL U781 ( .A(n686), .B(n678), .CI(n671), .CO(n352), .S(n353) );
  CNIVX2 U782 ( .A(n763), .Z(n994) );
  CNR2XL U783 ( .A(n36), .B(n46), .Z(n862) );
  CNR2XL U784 ( .A(n36), .B(n50), .Z(n847) );
  CNR2XL U785 ( .A(n36), .B(n40), .Z(n877) );
  COR2XL U786 ( .A(n32), .B(n36), .Z(n1003) );
  CNR2XL U787 ( .A(n36), .B(n52), .Z(n838) );
  CNR2XL U788 ( .A(n36), .B(n48), .Z(n855) );
  CNR2XL U789 ( .A(n36), .B(n28), .Z(n649) );
  CNR2XL U790 ( .A(n36), .B(n911), .Z(n805) );
  CNR2XL U791 ( .A(n36), .B(n27), .Z(n653) );
  CNR2XL U792 ( .A(n34), .B(n36), .Z(n883) );
  CNR2XL U793 ( .A(n36), .B(n24), .Z(n671) );
  CNR2XL U794 ( .A(n36), .B(n15), .Z(n778) );
  CNR2XL U795 ( .A(n36), .B(n16), .Z(n763) );
  COND1X2 U796 ( .A(n102), .B(n104), .C(n103), .Z(n101) );
  CANR1X2 U797 ( .A(n105), .B(n113), .C(n106), .Z(n104) );
  CANR1X2 U798 ( .A(n202), .B(n1007), .C(n199), .Z(n197) );
  COND1X1 U799 ( .A(n203), .B(n205), .C(n204), .Z(n202) );
  CIVXL U800 ( .A(n181), .Z(n180) );
  CANR1X1 U801 ( .A(n1000), .B(n186), .C(n183), .Z(n181) );
  COND1X1 U802 ( .A(n114), .B(n126), .C(n115), .Z(n113) );
  CANR1X1 U803 ( .A(n146), .B(n127), .C(n128), .Z(n126) );
  CNR2XL U804 ( .A(n40), .B(n24), .Z(n669) );
  CNR2XL U805 ( .A(n52), .B(n18), .Z(n726) );
  CNR2XL U806 ( .A(n50), .B(n19), .Z(n714) );
  CNR2XL U807 ( .A(n36), .B(n25), .Z(n664) );
  CNR2XL U808 ( .A(n34), .B(n17), .Z(n749) );
  CNR2XL U809 ( .A(n42), .B(n25), .Z(n661) );
  CNR2XL U810 ( .A(n40), .B(n22), .Z(n686) );
  CNR2XL U811 ( .A(n910), .B(n15), .Z(n766) );
  CNR2X1 U812 ( .A(n38), .B(n40), .Z(n876) );
  CNR2X1 U813 ( .A(n38), .B(n16), .Z(n762) );
  CNR2XL U814 ( .A(n32), .B(n40), .Z(n879) );
  CNR2XL U815 ( .A(n48), .B(n16), .Z(n757) );
  CNR2XL U816 ( .A(n48), .B(n54), .Z(n822) );
  CND2XL U817 ( .A(n1058), .B(n225), .Z(n132) );
  CEOXL U818 ( .A(n197), .B(n80), .Z(product[7]) );
  CANR1XL U819 ( .A(n210), .B(n1004), .C(n207), .Z(n205) );
  CNR2XL U820 ( .A(n42), .B(n15), .Z(n775) );
  CNR2XL U821 ( .A(n38), .B(n912), .Z(n816) );
  CNR2XL U822 ( .A(n40), .B(n52), .Z(n836) );
  CNR2XL U823 ( .A(n50), .B(n42), .Z(n844) );
  CNR2XL U824 ( .A(n36), .B(n912), .Z(n817) );
  CNR2X1 U825 ( .A(n34), .B(n23), .Z(n680) );
  CNR2XL U826 ( .A(n32), .B(n52), .Z(n840) );
  CNR2XL U827 ( .A(n46), .B(n42), .Z(n859) );
  CNR2XL U828 ( .A(n38), .B(n44), .Z(n867) );
  CNR2XL U829 ( .A(n40), .B(n912), .Z(n815) );
  CNR2XL U830 ( .A(n32), .B(n28), .Z(n651) );
  CNR2XL U831 ( .A(n36), .B(n44), .Z(n868) );
  CNR2XL U832 ( .A(n911), .B(n52), .Z(n797) );
  CNR2XL U833 ( .A(n46), .B(n52), .Z(n833) );
  CNR2XL U834 ( .A(n44), .B(n42), .Z(n865) );
  CNR2XL U835 ( .A(n42), .B(n52), .Z(n835) );
  CNR2XL U836 ( .A(n32), .B(n44), .Z(n870) );
  CNR2XL U837 ( .A(n32), .B(n30), .Z(n646) );
  CNR2XL U838 ( .A(n36), .B(n38), .Z(n880) );
  CIVX2 U839 ( .A(b[13]), .Z(n911) );
  CIVX2 U840 ( .A(b[15]), .Z(n15) );
  CIVX3 U841 ( .A(b[9]), .Z(n50) );
  CND2XL U842 ( .A(n885), .B(a[1]), .Z(n213) );
  CND2XL U843 ( .A(n1000), .B(n185), .Z(n77) );
  CNR2XL U844 ( .A(n427), .B(n446), .Z(n107) );
  CNR2XL U845 ( .A(n447), .B(n466), .Z(n110) );
  CNR2XL U846 ( .A(n467), .B(n484), .Z(n118) );
  CNR2XL U847 ( .A(n162), .B(n165), .Z(n160) );
  CNR2XL U848 ( .A(n503), .B(n518), .Z(n129) );
  CNR2XL U849 ( .A(n535), .B(n548), .Z(n139) );
  CND2XL U850 ( .A(n485), .B(n502), .Z(n124) );
  CND2XL U851 ( .A(n503), .B(n518), .Z(n130) );
  CND2XL U852 ( .A(n999), .B(n174), .Z(n75) );
  CND2XL U853 ( .A(n535), .B(n548), .Z(n140) );
  CND2XL U854 ( .A(n998), .B(n179), .Z(n76) );
  CND2XL U855 ( .A(n549), .B(n562), .Z(n152) );
  CND2XL U856 ( .A(n519), .B(n534), .Z(n137) );
  CND2IXL U857 ( .B(n162), .A(n163), .Z(n73) );
  CIVXL U858 ( .A(n179), .Z(n177) );
  CND2XL U859 ( .A(n233), .B(n188), .Z(n78) );
  CND2XL U860 ( .A(n235), .B(n196), .Z(n80) );
  CND2XL U861 ( .A(n1002), .B(n193), .Z(n79) );
  CND2XL U862 ( .A(n575), .B(n586), .Z(n163) );
  CND2XL U863 ( .A(n563), .B(n574), .Z(n157) );
  CND2XL U864 ( .A(n237), .B(n204), .Z(n82) );
  CND2XL U865 ( .A(n1004), .B(n209), .Z(n83) );
  CND2XL U866 ( .A(n1007), .B(n201), .Z(n81) );
  CNR2XL U867 ( .A(n34), .B(n44), .Z(n869) );
  CNR2XL U868 ( .A(n36), .B(n910), .Z(n792) );
  CNR2XL U869 ( .A(n34), .B(n28), .Z(n650) );
  CNR2XL U870 ( .A(n911), .B(n16), .Z(n752) );
  CNR2XL U871 ( .A(n44), .B(n21), .Z(n694) );
  CNR2XL U872 ( .A(n50), .B(n18), .Z(n727) );
  CNR2XL U873 ( .A(n46), .B(n23), .Z(n674) );
  CNR2XL U874 ( .A(n38), .B(n27), .Z(n652) );
  CNR2XL U875 ( .A(n50), .B(n21), .Z(n691) );
  CNR2XL U876 ( .A(n40), .B(n26), .Z(n656) );
  CNR2XL U877 ( .A(n54), .B(n19), .Z(n712) );
  CNR2XL U878 ( .A(n34), .B(n50), .Z(n848) );
  CNR2XL U879 ( .A(n32), .B(n27), .Z(n655) );
  CNR2XL U880 ( .A(n54), .B(n16), .Z(n754) );
  CNR2XL U881 ( .A(n42), .B(n22), .Z(n685) );
  CNR2XL U882 ( .A(n40), .B(n54), .Z(n826) );
  CNR2XL U883 ( .A(n46), .B(n21), .Z(n693) );
  CNR2XL U884 ( .A(n38), .B(n22), .Z(n687) );
  CNR2XL U885 ( .A(n44), .B(n19), .Z(n717) );
  CEOXL U886 ( .A(n213), .B(n1003), .Z(product[3]) );
  CNR2XL U887 ( .A(n38), .B(n17), .Z(n747) );
  CNR2XL U888 ( .A(n38), .B(n910), .Z(n791) );
  CNR2XL U889 ( .A(n44), .B(n54), .Z(n824) );
  CNR2XL U890 ( .A(n38), .B(n54), .Z(n827) );
  CNR2XL U891 ( .A(n48), .B(n21), .Z(n692) );
  CNR2XL U892 ( .A(n52), .B(n19), .Z(n713) );
  CNR2XL U893 ( .A(n911), .B(n910), .Z(n781) );
  CNR2XL U894 ( .A(n36), .B(n22), .Z(n688) );
  CNR2XL U895 ( .A(n38), .B(n21), .Z(n697) );
  CNR2XL U896 ( .A(n44), .B(n17), .Z(n744) );
  CNR2XL U897 ( .A(n50), .B(n910), .Z(n785) );
  CNR2XL U898 ( .A(n54), .B(n912), .Z(n808) );
  CNR2XL U899 ( .A(n42), .B(n20), .Z(n706) );
  CNR2XL U900 ( .A(n54), .B(n910), .Z(n783) );
  CNR2XL U901 ( .A(n46), .B(n19), .Z(n716) );
  CNR2XL U902 ( .A(n46), .B(n18), .Z(n729) );
  CNR2XL U903 ( .A(n48), .B(n17), .Z(n742) );
  CNR2XL U904 ( .A(n50), .B(n16), .Z(n756) );
  CNR2XL U905 ( .A(n50), .B(n54), .Z(n821) );
  CNR2XL U906 ( .A(n34), .B(n25), .Z(n665) );
  CNR2XL U907 ( .A(n912), .B(n910), .Z(n782) );
  CNR2XL U908 ( .A(n32), .B(n910), .Z(n794) );
  CNR2XL U909 ( .A(n46), .B(n54), .Z(n823) );
  CNR2XL U910 ( .A(n34), .B(n911), .Z(n806) );
  CNR2XL U911 ( .A(n38), .B(n26), .Z(n657) );
  CNR2XL U912 ( .A(n46), .B(n22), .Z(n683) );
  CNR2XL U913 ( .A(n54), .B(n18), .Z(n725) );
  CNR2XL U914 ( .A(n34), .B(n48), .Z(n856) );
  CNR2XL U915 ( .A(n54), .B(n17), .Z(n739) );
  CNR2XL U916 ( .A(n42), .B(n18), .Z(n731) );
  CNR2XL U917 ( .A(n40), .B(n19), .Z(n719) );
  CNR2XL U918 ( .A(n34), .B(n912), .Z(n818) );
  CNR2XL U919 ( .A(n36), .B(n54), .Z(n828) );
  CNR2XL U920 ( .A(n42), .B(n19), .Z(n718) );
  CNR2XL U921 ( .A(n34), .B(n22), .Z(n689) );
  CNR2XL U922 ( .A(n46), .B(n16), .Z(n758) );
  CNR2XL U923 ( .A(n52), .B(n17), .Z(n740) );
  CNR2XL U924 ( .A(n34), .B(n26), .Z(n659) );
  CNR2XL U925 ( .A(n911), .B(n17), .Z(n737) );
  CNR2XL U926 ( .A(n44), .B(n24), .Z(n667) );
  CNR2XL U927 ( .A(n52), .B(n20), .Z(n701) );
  CNR2XL U928 ( .A(n32), .B(n34), .Z(n885) );
  CNR2XL U929 ( .A(n40), .B(n17), .Z(n746) );
  CNR2XL U930 ( .A(n48), .B(n19), .Z(n715) );
  CNR2XL U931 ( .A(n34), .B(n54), .Z(n829) );
  CNR2XL U932 ( .A(n34), .B(n24), .Z(n672) );
  CNR2XL U933 ( .A(n36), .B(n23), .Z(n679) );
  CNR2XL U934 ( .A(n40), .B(n21), .Z(n696) );
  CNR2XL U935 ( .A(n34), .B(n38), .Z(n881) );
  CNR2XL U936 ( .A(n34), .B(n15), .Z(n779) );
  CNR2XL U937 ( .A(n36), .B(n20), .Z(n709) );
  CNR2XL U938 ( .A(n38), .B(n25), .Z(n663) );
  CNR2XL U939 ( .A(n34), .B(n46), .Z(n863) );
  CNR2XL U940 ( .A(n34), .B(n16), .Z(n764) );
  CNR2XL U941 ( .A(n46), .B(n17), .Z(n743) );
  CNR2XL U942 ( .A(n32), .B(n54), .Z(n830) );
  CNR2XL U943 ( .A(n44), .B(n18), .Z(n730) );
  CNR2XL U944 ( .A(n910), .B(n52), .Z(n784) );
  CNR2XL U945 ( .A(n36), .B(n21), .Z(n698) );
  CNR2XL U946 ( .A(n34), .B(n910), .Z(n793) );
  CNR2XL U947 ( .A(n50), .B(n17), .Z(n741) );
  CNR2XL U948 ( .A(n48), .B(n18), .Z(n728) );
  CNR2XL U949 ( .A(n34), .B(n42), .Z(n874) );
  CNR2XL U950 ( .A(n32), .B(n18), .Z(n736) );
  CNR2XL U951 ( .A(n40), .B(n910), .Z(n790) );
  CNR2XL U952 ( .A(n34), .B(n29), .Z(n647) );
  CNR2XL U953 ( .A(n912), .B(n18), .Z(n724) );
  CEO3X1 U954 ( .A(n724), .B(n280), .C(n278), .Z(n248) );
  CNR2XL U955 ( .A(n912), .B(n17), .Z(n738) );
  CNR2XL U956 ( .A(n910), .B(n16), .Z(n751) );
  CEO3X1 U957 ( .A(n661), .B(n652), .C(n656), .Z(n251) );
  CNR2XL U958 ( .A(n48), .B(n22), .Z(n682) );
  CEO3X1 U959 ( .A(n737), .B(n691), .C(n712), .Z(n249) );
  CNR2XL U960 ( .A(n34), .B(n40), .Z(n878) );
  CIVX4 U961 ( .A(b[3]), .Z(n38) );
  CIVX4 U962 ( .A(b[4]), .Z(n40) );
  CNR2XL U963 ( .A(n132), .B(n1045), .Z(n127) );
  CIVX4 U964 ( .A(b[6]), .Z(n44) );
  CIVX4 U965 ( .A(b[5]), .Z(n42) );
  CIVX4 U966 ( .A(b[7]), .Z(n46) );
  CIVX4 U967 ( .A(b[8]), .Z(n48) );
  CIVX4 U968 ( .A(b[10]), .Z(n52) );
  CIVX3 U969 ( .A(b[12]), .Z(n912) );
  CNR2XL U970 ( .A(n40), .B(n42), .Z(n871) );
  CIVX1 U971 ( .A(b[28]), .Z(n28) );
  CIVXL U972 ( .A(n1043), .Z(n135) );
  CND2IXL U973 ( .B(n212), .A(n213), .Z(n84) );
  CENX1 U974 ( .A(n77), .B(n186), .Z(product[10]) );
  COND1XL U975 ( .A(n181), .B(n169), .C(n170), .Z(n168) );
  CND2X1 U976 ( .A(n999), .B(n998), .Z(n169) );
  CANR1XL U977 ( .A(n177), .B(n999), .C(n172), .Z(n170) );
  COND1XL U978 ( .A(n166), .B(n162), .C(n163), .Z(n161) );
  COR2X1 U979 ( .A(n549), .B(n562), .Z(n995) );
  CND2XL U980 ( .A(n427), .B(n446), .Z(n108) );
  CND2XL U981 ( .A(n467), .B(n484), .Z(n119) );
  CND2XL U982 ( .A(n447), .B(n466), .Z(n111) );
  COR2X1 U983 ( .A(n519), .B(n534), .Z(n996) );
  COR2X1 U984 ( .A(n485), .B(n502), .Z(n997) );
  CANR1XL U985 ( .A(n194), .B(n1002), .C(n191), .Z(n189) );
  COND1XL U986 ( .A(n195), .B(n197), .C(n196), .Z(n194) );
  COND1XL U987 ( .A(n187), .B(n189), .C(n188), .Z(n186) );
  CNR2X1 U988 ( .A(n575), .B(n586), .Z(n162) );
  CENX1 U989 ( .A(n79), .B(n194), .Z(product[8]) );
  CNR2X1 U990 ( .A(n587), .B(n596), .Z(n165) );
  CEOXL U991 ( .A(n189), .B(n78), .Z(product[9]) );
  COR2X1 U992 ( .A(n607), .B(n614), .Z(n998) );
  COR2X1 U993 ( .A(n597), .B(n606), .Z(n999) );
  CND2X1 U994 ( .A(n597), .B(n606), .Z(n174) );
  CND2X1 U995 ( .A(n615), .B(n622), .Z(n185) );
  CND2X1 U996 ( .A(n607), .B(n614), .Z(n179) );
  COR2X1 U997 ( .A(n615), .B(n622), .Z(n1000) );
  CND2X1 U998 ( .A(n587), .B(n596), .Z(n166) );
  COR2X1 U999 ( .A(n563), .B(n574), .Z(n1001) );
  CENX1 U1000 ( .A(n81), .B(n202), .Z(product[6]) );
  CND2X1 U1001 ( .A(n1006), .B(n92), .Z(n60) );
  CNR2X1 U1002 ( .A(n635), .B(n638), .Z(n195) );
  CNR2X1 U1003 ( .A(n623), .B(n628), .Z(n187) );
  CEOXL U1004 ( .A(n205), .B(n82), .Z(product[5]) );
  CND2X1 U1005 ( .A(n629), .B(n634), .Z(n193) );
  CND2X1 U1006 ( .A(n635), .B(n638), .Z(n196) );
  CND2X1 U1007 ( .A(n623), .B(n628), .Z(n188) );
  COR2X1 U1008 ( .A(n629), .B(n634), .Z(n1002) );
  CENX1 U1009 ( .A(n83), .B(n210), .Z(product[4]) );
  CNR2X1 U1010 ( .A(n213), .B(n1003), .Z(n210) );
  CNR2X1 U1011 ( .A(n32), .B(n38), .Z(n882) );
  CNR2X1 U1012 ( .A(n40), .B(n46), .Z(n860) );
  CNR2X1 U1013 ( .A(n42), .B(n24), .Z(n668) );
  CNR2X1 U1014 ( .A(n40), .B(n48), .Z(n853) );
  CNR2X1 U1015 ( .A(n48), .B(n911), .Z(n799) );
  CNR2X1 U1016 ( .A(n50), .B(n912), .Z(n810) );
  CNR2X1 U1017 ( .A(n54), .B(n52), .Z(n820) );
  CNR2X1 U1018 ( .A(n38), .B(n911), .Z(n804) );
  CNR2X1 U1019 ( .A(n32), .B(n16), .Z(n765) );
  CNR2X1 U1020 ( .A(n54), .B(n42), .Z(n825) );
  CNR2X1 U1021 ( .A(n912), .B(n15), .Z(n768) );
  CNR2X1 U1022 ( .A(n40), .B(n23), .Z(n677) );
  CENX1 U1023 ( .A(n101), .B(n62), .Z(product[25]) );
  CND2X1 U1024 ( .A(n1009), .B(n100), .Z(n62) );
  CNR2X1 U1025 ( .A(n911), .B(n42), .Z(n802) );
  CNR2X1 U1026 ( .A(n48), .B(n50), .Z(n841) );
  CNR2X1 U1027 ( .A(n40), .B(n911), .Z(n803) );
  CNR2X1 U1028 ( .A(n912), .B(n42), .Z(n814) );
  CNR2X1 U1029 ( .A(n46), .B(n910), .Z(n787) );
  CNR2X1 U1030 ( .A(n44), .B(n15), .Z(n774) );
  CNR2X1 U1031 ( .A(n38), .B(n18), .Z(n733) );
  CNR2X1 U1032 ( .A(n42), .B(n23), .Z(n676) );
  CNR2X1 U1033 ( .A(n46), .B(n48), .Z(n850) );
  CNR2X1 U1034 ( .A(n52), .B(n15), .Z(n770) );
  CNR2X1 U1035 ( .A(n44), .B(n48), .Z(n851) );
  CNR2X1 U1036 ( .A(n643), .B(n644), .Z(n203) );
  CNR2X1 U1037 ( .A(n36), .B(n19), .Z(n721) );
  CNR2X1 U1038 ( .A(n42), .B(n16), .Z(n760) );
  CNR2X1 U1039 ( .A(n32), .B(n21), .Z(n700) );
  CNR2X1 U1040 ( .A(n48), .B(n52), .Z(n832) );
  CNR2X1 U1041 ( .A(n44), .B(n911), .Z(n801) );
  CNR2X1 U1042 ( .A(n46), .B(n912), .Z(n812) );
  CNR2X1 U1043 ( .A(n50), .B(n52), .Z(n831) );
  CNR2X1 U1044 ( .A(n46), .B(n50), .Z(n842) );
  CNR2X1 U1045 ( .A(n44), .B(n52), .Z(n834) );
  CNR2X1 U1046 ( .A(n44), .B(n46), .Z(n858) );
  CNR2X1 U1047 ( .A(n32), .B(n911), .Z(n807) );
  CNR2X1 U1048 ( .A(n38), .B(n52), .Z(n837) );
  CNR2X1 U1049 ( .A(n912), .B(n911), .Z(n795) );
  CNR2X1 U1050 ( .A(n52), .B(n16), .Z(n755) );
  CNR2X1 U1051 ( .A(n42), .B(n21), .Z(n695) );
  CNR2X1 U1052 ( .A(n48), .B(n910), .Z(n786) );
  CNR2X1 U1053 ( .A(n912), .B(n52), .Z(n809) );
  CNR2X1 U1054 ( .A(n40), .B(n18), .Z(n732) );
  CNR2X1 U1055 ( .A(n40), .B(n44), .Z(n866) );
  CNR2X1 U1056 ( .A(n38), .B(n46), .Z(n861) );
  CNR2X1 U1057 ( .A(n38), .B(n48), .Z(n854) );
  CNR2X1 U1058 ( .A(n911), .B(n15), .Z(n767) );
  CNR2X1 U1059 ( .A(n48), .B(n20), .Z(n703) );
  CNR2X1 U1060 ( .A(n34), .B(n27), .Z(n654) );
  CNR2X1 U1061 ( .A(n38), .B(n19), .Z(n720) );
  CNR2X1 U1062 ( .A(n32), .B(n22), .Z(n690) );
  CNR2X1 U1063 ( .A(n34), .B(n21), .Z(n699) );
  CNR2X1 U1064 ( .A(n32), .B(n48), .Z(n857) );
  CNR2X1 U1065 ( .A(n38), .B(n42), .Z(n872) );
  CEOXL U1066 ( .A(n61), .B(n96), .Z(product[26]) );
  CND2X1 U1067 ( .A(n216), .B(n95), .Z(n61) );
  CNR2X1 U1068 ( .A(n912), .B(n16), .Z(n753) );
  CNR2X1 U1069 ( .A(n44), .B(n22), .Z(n684) );
  CNR2X1 U1070 ( .A(n32), .B(n23), .Z(n681) );
  CNR2X1 U1071 ( .A(n48), .B(n912), .Z(n811) );
  CNR2X1 U1072 ( .A(n36), .B(n18), .Z(n734) );
  CNR2X1 U1073 ( .A(n34), .B(n19), .Z(n722) );
  CNR2X1 U1074 ( .A(n32), .B(n24), .Z(n673) );
  CNR2X1 U1075 ( .A(n44), .B(n50), .Z(n843) );
  CNR2X1 U1076 ( .A(n40), .B(n15), .Z(n776) );
  CNR2X1 U1077 ( .A(n36), .B(n17), .Z(n748) );
  CNR2X1 U1078 ( .A(n910), .B(n42), .Z(n789) );
  COR2X1 U1079 ( .A(n645), .B(n882), .Z(n1004) );
  CNR2X1 U1080 ( .A(n50), .B(n911), .Z(n798) );
  CAOR1X1 U1081 ( .A(n1006), .B(n93), .C(n90), .Z(n1005) );
  CNR2X1 U1082 ( .A(n38), .B(n24), .Z(n670) );
  CNR2X1 U1083 ( .A(n44), .B(n912), .Z(n813) );
  CNR2X1 U1084 ( .A(n38), .B(n15), .Z(n777) );
  CNR2X1 U1085 ( .A(n40), .B(n50), .Z(n845) );
  CNR2X1 U1086 ( .A(n38), .B(n23), .Z(n678) );
  CNR2X1 U1087 ( .A(n32), .B(n19), .Z(n723) );
  CNR2X1 U1088 ( .A(n32), .B(n50), .Z(n849) );
  CNR2X1 U1089 ( .A(n38), .B(n50), .Z(n846) );
  CNR2X1 U1090 ( .A(n32), .B(n46), .Z(n864) );
  CNR2X1 U1091 ( .A(n48), .B(n15), .Z(n772) );
  CNR2X1 U1092 ( .A(n54), .B(n15), .Z(n769) );
  CNR2X1 U1093 ( .A(n32), .B(n26), .Z(n660) );
  CNR2X1 U1094 ( .A(n44), .B(n20), .Z(n705) );
  CNR2X1 U1095 ( .A(n46), .B(n911), .Z(n800) );
  CNR2X1 U1096 ( .A(n44), .B(n910), .Z(n788) );
  CNR2X1 U1097 ( .A(n40), .B(n16), .Z(n761) );
  CNR2X1 U1098 ( .A(n50), .B(n20), .Z(n702) );
  CNR2X1 U1099 ( .A(n32), .B(n29), .Z(n648) );
  CNR2X1 U1100 ( .A(n50), .B(n15), .Z(n771) );
  CNR2X1 U1101 ( .A(n44), .B(n16), .Z(n759) );
  CNR2X1 U1102 ( .A(n46), .B(n15), .Z(n773) );
  CNR2X1 U1103 ( .A(n42), .B(n17), .Z(n745) );
  CNR2X1 U1104 ( .A(n54), .B(n911), .Z(n796) );
  CNR2X1 U1105 ( .A(n40), .B(n20), .Z(n707) );
  CNR2X1 U1106 ( .A(n32), .B(n912), .Z(n819) );
  CEOX1 U1107 ( .A(n646), .B(n647), .Z(n253) );
  CND2X1 U1108 ( .A(n645), .B(n882), .Z(n209) );
  CND2X1 U1109 ( .A(n639), .B(n641), .Z(n201) );
  CND2X1 U1110 ( .A(n335), .B(n358), .Z(n92) );
  CNR2X1 U1111 ( .A(n44), .B(n23), .Z(n675) );
  CND2X1 U1112 ( .A(n643), .B(n644), .Z(n204) );
  COR2X1 U1113 ( .A(n335), .B(n358), .Z(n1006) );
  COR2X1 U1114 ( .A(n639), .B(n641), .Z(n1007) );
  CEOXL U1115 ( .A(n63), .B(n104), .Z(product[24]) );
  CND2X1 U1116 ( .A(n218), .B(n103), .Z(n63) );
  CNR2XL U1117 ( .A(n1052), .B(n1050), .Z(n105) );
  COND1XL U1118 ( .A(n1049), .B(n1052), .C(n1051), .Z(n106) );
  COND1XL U1119 ( .A(n1045), .B(n133), .C(n1044), .Z(n128) );
  CIVX4 U1120 ( .A(b[1]), .Z(n34) );
  CND2XL U1121 ( .A(n1057), .B(n1056), .Z(n147) );
  CND2XL U1122 ( .A(n221), .B(n1059), .Z(n114) );
  CANR1XL U1123 ( .A(n122), .B(n221), .C(n117), .Z(n115) );
  CANR1XL U1124 ( .A(n142), .B(n1058), .C(n135), .Z(n133) );
  CIVX2 U1125 ( .A(b[21]), .Z(n21) );
  CIVX2 U1126 ( .A(b[11]), .Z(n54) );
  CIVX2 U1127 ( .A(b[22]), .Z(n22) );
  CIVX2 U1128 ( .A(b[14]), .Z(n910) );
  CIVX2 U1129 ( .A(b[16]), .Z(n16) );
  CNR2X1 U1130 ( .A(n1011), .B(n1010), .Z(n102) );
  CNR2X1 U1131 ( .A(n359), .B(n1015), .Z(n94) );
  CIVX2 U1132 ( .A(b[18]), .Z(n18) );
  CNR2XL U1133 ( .A(n38), .B(n20), .Z(n708) );
  CNR2XL U1134 ( .A(n32), .B(n42), .Z(n875) );
  CNR2XL U1135 ( .A(n34), .B(n52), .Z(n839) );
  CENX1 U1136 ( .A(n1008), .B(n85), .Z(product[31]) );
  CENX1 U1137 ( .A(n1030), .B(n254), .Z(n1008) );
  CIVX2 U1138 ( .A(b[19]), .Z(n19) );
  CIVX2 U1139 ( .A(b[20]), .Z(n20) );
  COR2X1 U1140 ( .A(n1014), .B(n1012), .Z(n1009) );
  CNR2X1 U1141 ( .A(n34), .B(n20), .Z(n710) );
  CNR2XL U1142 ( .A(n40), .B(n25), .Z(n662) );
  CNR2X1 U1143 ( .A(n46), .B(n20), .Z(n704) );
  CNR2XL U1144 ( .A(n34), .B(n18), .Z(n735) );
  CNR2XL U1145 ( .A(n48), .B(n42), .Z(n852) );
  CNR2XL U1146 ( .A(n32), .B(n25), .Z(n666) );
  CNR2XL U1147 ( .A(n36), .B(n42), .Z(n873) );
  CNR2XL U1148 ( .A(n32), .B(n15), .Z(n780) );
  CND2X1 U1149 ( .A(n1014), .B(n1012), .Z(n100) );
  CND2X1 U1150 ( .A(n1011), .B(n1010), .Z(n103) );
  CND2X1 U1151 ( .A(n359), .B(n1015), .Z(n95) );
  CEOX1 U1152 ( .A(n71), .B(n153), .Z(product[16]) );
  CND2XL U1153 ( .A(n1057), .B(n1040), .Z(n71) );
  CANR1XL U1154 ( .A(n1056), .B(n158), .C(n155), .Z(n153) );
  CENX1 U1155 ( .A(n138), .B(n69), .Z(product[18]) );
  CND2XL U1156 ( .A(n1058), .B(n1043), .Z(n69) );
  COND1XL U1157 ( .A(n1042), .B(n145), .C(n1041), .Z(n138) );
  CENX1 U1158 ( .A(n131), .B(n68), .Z(product[19]) );
  CND2XL U1159 ( .A(n223), .B(n1044), .Z(n68) );
  COND1XL U1160 ( .A(n132), .B(n145), .C(n133), .Z(n131) );
  CENX1 U1161 ( .A(n109), .B(n64), .Z(product[23]) );
  CND2XL U1162 ( .A(n219), .B(n1051), .Z(n64) );
  COND1XL U1163 ( .A(n1050), .B(n112), .C(n1049), .Z(n109) );
  CENX1 U1164 ( .A(n1033), .B(n1053), .Z(n1094) );
  CENX1 U1165 ( .A(n164), .B(n1037), .Z(n1091) );
  COND1XL U1166 ( .A(n1036), .B(n167), .C(n1035), .Z(n164) );
  CENX1 U1167 ( .A(n158), .B(n72), .Z(product[15]) );
  CND2XL U1168 ( .A(n1056), .B(n1039), .Z(n72) );
  CENX1 U1169 ( .A(n125), .B(n67), .Z(product[20]) );
  CND2XL U1170 ( .A(n1059), .B(n1046), .Z(n67) );
  CEOX1 U1171 ( .A(n175), .B(n1034), .Z(n1093) );
  CANR1XL U1172 ( .A(n1055), .B(n1053), .C(n1054), .Z(n175) );
  CEOX1 U1173 ( .A(n74), .B(n167), .Z(n1092) );
  CND2X1 U1174 ( .A(n229), .B(n1035), .Z(n74) );
  CEOX1 U1175 ( .A(n70), .B(n145), .Z(product[17]) );
  CND2XL U1176 ( .A(n225), .B(n1041), .Z(n70) );
  CEOX1 U1177 ( .A(n66), .B(n120), .Z(product[21]) );
  CND2XL U1178 ( .A(n221), .B(n1047), .Z(n66) );
  CANR1XL U1179 ( .A(n1059), .B(n125), .C(n122), .Z(n120) );
  CEOX1 U1180 ( .A(n65), .B(n112), .Z(product[22]) );
  CNR2XL U1181 ( .A(n885), .B(a[1]), .Z(n212) );
  CIVX2 U1182 ( .A(n84), .Z(product[2]) );
  CIVX2 U1183 ( .A(n100), .Z(n98) );
  CIVX2 U1184 ( .A(n92), .Z(n90) );
  CIVX2 U1185 ( .A(b[30]), .Z(n30) );
  CIVX2 U1186 ( .A(b[29]), .Z(n29) );
  CIVX2 U1187 ( .A(b[27]), .Z(n27) );
  CIVX2 U1188 ( .A(b[26]), .Z(n26) );
  CIVX2 U1189 ( .A(b[25]), .Z(n25) );
  CIVX2 U1190 ( .A(b[24]), .Z(n24) );
  CIVX2 U1191 ( .A(n203), .Z(n237) );
  CIVX2 U1192 ( .A(n195), .Z(n235) );
  CIVX2 U1193 ( .A(n187), .Z(n233) );
  CIVX2 U1194 ( .A(b[23]), .Z(n23) );
  CIVX2 U1195 ( .A(n1036), .Z(n229) );
  CIVX2 U1196 ( .A(n1045), .Z(n223) );
  CIVX2 U1197 ( .A(n1050), .Z(n220) );
  CIVX2 U1198 ( .A(n1052), .Z(n219) );
  CIVX2 U1199 ( .A(n102), .Z(n218) );
  CIVX2 U1200 ( .A(n94), .Z(n216) );
  CIVX2 U1201 ( .A(n209), .Z(n207) );
  CIVX2 U1202 ( .A(n201), .Z(n199) );
  CIVX2 U1203 ( .A(n193), .Z(n191) );
  CIVX2 U1204 ( .A(n185), .Z(n183) );
  CIVX2 U1205 ( .A(n174), .Z(n172) );
  CIVX2 U1206 ( .A(n1031), .Z(n167) );
  CIVX2 U1207 ( .A(n1039), .Z(n155) );
  CIVX2 U1208 ( .A(n1040), .Z(n150) );
  CIVX2 U1209 ( .A(n146), .Z(n145) );
  CIVX2 U1210 ( .A(n1041), .Z(n142) );
  CIVX2 U1211 ( .A(n1042), .Z(n225) );
  CIVX2 U1212 ( .A(n126), .Z(n125) );
  CIVX2 U1213 ( .A(n1046), .Z(n122) );
  CIVX2 U1214 ( .A(n1047), .Z(n117) );
  CIVX2 U1215 ( .A(n1048), .Z(n221) );
endmodule


module calc_DW02_mult_2_stage_8 ( A, B, TC, CLK, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC, CLK;
  wire   n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, \B_extended[32] ,
         n6, n8, n10, n12, n14, n16, n18, n20, n22, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34;
  assign \B_extended[32]  = B[31];

  calc_DW_mult_tc_19 mult_96 ( .a({\B_extended[32] , A}), .b({\B_extended[32] , 
        \B_extended[32] , B[30:0]}), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, PRODUCT[31:11], n35, n36, n37, n38, n39, n40, 
        n41, n42, n43, SYNOPSYS_UNCONNECTED__34, n44}), .dw3_CLK(CLK) );
  CFD1QXL clk_r_REG56_S1 ( .D(n43), .CP(CLK), .Q(n26) );
  CFD1QXL clk_r_REG57_S1 ( .D(n42), .CP(CLK), .Q(n27) );
  CFD1QXL clk_r_REG52_S1 ( .D(n39), .CP(CLK), .Q(n30) );
  CFD1QXL clk_r_REG55_S1 ( .D(n40), .CP(CLK), .Q(n29) );
  CFD1QXL clk_r_REG54_S1 ( .D(n41), .CP(CLK), .Q(n28) );
  CFD1QXL clk_r_REG51_S1 ( .D(n36), .CP(CLK), .Q(n33) );
  CFD1QXL clk_r_REG50_S1 ( .D(n37), .CP(CLK), .Q(n32) );
  CFD1QXL clk_r_REG53_S1 ( .D(n38), .CP(CLK), .Q(n31) );
  CFD1QXL clk_r_REG45_S1 ( .D(n35), .CP(CLK), .Q(n34) );
  CFD1QXL clk_r_REG59_S1 ( .D(n44), .CP(CLK), .Q(n25) );
  CIVDXL U1 ( .A(n30), .Z1(n6) );
  CNIVX1 U2 ( .A(n6), .Z(PRODUCT[6]) );
  CIVDXL U3 ( .A(n25), .Z1(n8) );
  CNIVX1 U4 ( .A(n8), .Z(PRODUCT[0]) );
  CIVDXL U5 ( .A(n28), .Z1(n10) );
  CNIVX1 U6 ( .A(n10), .Z(PRODUCT[4]) );
  CIVDXL U7 ( .A(n27), .Z1(n12) );
  CNIVX1 U8 ( .A(n12), .Z(PRODUCT[3]) );
  CIVDXL U9 ( .A(n26), .Z1(n14) );
  CNIVX1 U10 ( .A(n14), .Z(PRODUCT[2]) );
  CIVDXL U11 ( .A(n33), .Z1(n16) );
  CNIVX1 U12 ( .A(n16), .Z(PRODUCT[9]) );
  CIVDXL U13 ( .A(n32), .Z1(n18) );
  CNIVX1 U14 ( .A(n18), .Z(PRODUCT[8]) );
  CIVDXL U15 ( .A(n31), .Z1(n20) );
  CNIVX1 U16 ( .A(n20), .Z(PRODUCT[7]) );
  CIVDXL U17 ( .A(n29), .Z1(n22) );
  CNIVX1 U18 ( .A(n22), .Z(PRODUCT[5]) );
  CIVDXL U19 ( .A(n34), .Z1(n24) );
  CNIVX1 U20 ( .A(n24), .Z(PRODUCT[10]) );
endmodule


module calc_DW_mult_tc_20 ( a, b, product, dw2_CLK );
  input [32:0] a;
  input [32:0] b;
  output [65:0] product;
  input dw2_CLK;
  wire   n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n32, n34, n36, n38, n40, n42, n44, n46, n48, n50, n52, n54,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n90, n92, n93, n94, n95, n96, n98, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n117,
         n118, n119, n120, n122, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n135, n137, n138, n139, n140, n142, n145, n146,
         n147, n148, n150, n152, n153, n155, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n172, n174,
         n175, n177, n179, n180, n181, n183, n185, n186, n187, n188, n189,
         n191, n193, n194, n195, n196, n197, n199, n201, n202, n203, n204,
         n205, n207, n209, n210, n212, n213, n216, n218, n219, n220, n221,
         n223, n225, n229, n233, n235, n237, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n885, n910, n911, n912, \b[0] , n1091, n1090, n1089, n986, n987,
         n989, n991, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058;
  assign product[0] = \b[0] ;
  assign \b[0]  = b[0];
  assign n1058 = dw2_CLK;

  CFA1X1 U50 ( .A(n282), .B(n86), .CI(n255), .CO(n85), .S(product[30]) );
  CFA1X1 U51 ( .A(n308), .B(n87), .CI(n283), .CO(n86), .S(product[29]) );
  CFA1X1 U52 ( .A(n334), .B(n1004), .CI(n309), .CO(n87), .S(product[28]) );
  CEO3X2 U256 ( .A(n258), .B(n241), .C(n256), .Z(n240) );
  CEO3X2 U257 ( .A(n260), .B(n243), .C(n242), .Z(n241) );
  CEO3X2 U258 ( .A(n245), .B(n262), .C(n244), .Z(n242) );
  CEO3X2 U259 ( .A(n246), .B(n247), .C(n264), .Z(n243) );
  CEO3X2 U260 ( .A(n248), .B(n268), .C(n266), .Z(n244) );
  CEO3X2 U261 ( .A(n249), .B(n250), .C(n270), .Z(n245) );
  CEO3X2 U262 ( .A(n274), .B(n251), .C(n252), .Z(n246) );
  CEO3X2 U263 ( .A(n276), .B(n272), .C(n253), .Z(n247) );
  CEO3X2 U266 ( .A(n667), .B(n674), .C(n682), .Z(n250) );
  CEO3X2 U268 ( .A(n701), .B(n649), .C(n751), .Z(n252) );
  CFA1X1 U270 ( .A(n1026), .B(n1027), .CI(n1025), .CO(n254), .S(n255) );
  CFA1X1 U271 ( .A(n288), .B(n286), .CI(n261), .CO(n256), .S(n257) );
  CFA1X1 U272 ( .A(n265), .B(n263), .CI(n290), .CO(n258), .S(n259) );
  CFA1X1 U273 ( .A(n269), .B(n292), .CI(n267), .CO(n260), .S(n261) );
  CFA1X1 U274 ( .A(n271), .B(n294), .CI(n296), .CO(n262), .S(n263) );
  CFA1X1 U275 ( .A(n275), .B(n277), .CI(n273), .CO(n264), .S(n265) );
  CFA1X1 U276 ( .A(n298), .B(n279), .CI(n300), .CO(n266), .S(n267) );
  CFA1X1 U277 ( .A(n281), .B(n302), .CI(n304), .CO(n268), .S(n269) );
  CFA1X1 U278 ( .A(n692), .B(n306), .CI(n713), .CO(n270), .S(n271) );
  CFA1X1 U279 ( .A(n725), .B(n683), .CI(n657), .CO(n272), .S(n273) );
  CFA1X1 U280 ( .A(n668), .B(n653), .CI(n987), .CO(n274), .S(n275) );
  CFA1X1 U281 ( .A(n675), .B(n752), .CI(n650), .CO(n276), .S(n277) );
  CFA1X1 U282 ( .A(n702), .B(n766), .CI(n648), .CO(n278), .S(n279) );
  CHA1X1 U283 ( .A(a[15]), .B(n662), .CO(n280), .S(n281) );
  CFA1X1 U284 ( .A(n1023), .B(n1024), .CI(n1022), .CO(n282), .S(n283) );
  CFA1X1 U285 ( .A(n291), .B(n312), .CI(n289), .CO(n284), .S(n285) );
  CFA1X1 U286 ( .A(n316), .B(n314), .CI(n293), .CO(n286), .S(n287) );
  CFA1X1 U287 ( .A(n297), .B(n295), .CI(n318), .CO(n288), .S(n289) );
  CFA1X1 U288 ( .A(n301), .B(n320), .CI(n299), .CO(n290), .S(n291) );
  CFA1X1 U289 ( .A(n305), .B(n322), .CI(n303), .CO(n292), .S(n293) );
  CFA1X1 U290 ( .A(n328), .B(n326), .CI(n324), .CO(n294), .S(n295) );
  CFA1X1 U291 ( .A(n332), .B(n330), .CI(n307), .CO(n296), .S(n297) );
  CFA1X1 U292 ( .A(n714), .B(n693), .CI(n676), .CO(n298), .S(n299) );
  CFA1X1 U294 ( .A(n684), .B(n739), .CI(n753), .CO(n302), .S(n303) );
  CFA1X1 U295 ( .A(n703), .B(n654), .CI(n767), .CO(n304), .S(n305) );
  CHA1X1 U296 ( .A(n663), .B(n651), .CO(n306), .S(n307) );
  CFA1X1 U297 ( .A(n1020), .B(n1021), .CI(n1019), .CO(n308), .S(n309) );
  CFA1X1 U298 ( .A(n340), .B(n338), .CI(n315), .CO(n310), .S(n311) );
  CFA1X1 U299 ( .A(n342), .B(n317), .CI(n319), .CO(n312), .S(n313) );
  CFA1X1 U300 ( .A(n346), .B(n321), .CI(n344), .CO(n314), .S(n315) );
  CFA1X1 U301 ( .A(n331), .B(n323), .CI(n329), .CO(n316), .S(n317) );
  CFA1X1 U302 ( .A(n348), .B(n325), .CI(n327), .CO(n318), .S(n319) );
  CFA1X1 U303 ( .A(n354), .B(n352), .CI(n350), .CO(n320), .S(n321) );
  CFA1X1 U304 ( .A(n715), .B(n333), .CI(n356), .CO(n322), .S(n323) );
  CFA1X1 U305 ( .A(n727), .B(n694), .CI(n677), .CO(n324), .S(n325) );
  CFA1X1 U306 ( .A(n670), .B(n659), .CI(n740), .CO(n326), .S(n327) );
  CFA1X1 U307 ( .A(n685), .B(n754), .CI(n655), .CO(n328), .S(n329) );
  CFA1X1 U308 ( .A(n664), .B(n781), .CI(n768), .CO(n330), .S(n331) );
  CHA1X1 U309 ( .A(a[14]), .B(n704), .CO(n332), .S(n333) );
  CFA1X1 U310 ( .A(n1017), .B(n1018), .CI(n1016), .CO(n334), .S(n335) );
  CFA1X1 U311 ( .A(n364), .B(n362), .CI(n341), .CO(n336), .S(n337) );
  CFA1X1 U312 ( .A(n366), .B(n343), .CI(n345), .CO(n338), .S(n339) );
  CFA1X1 U313 ( .A(n370), .B(n347), .CI(n368), .CO(n340), .S(n341) );
  CFA1X1 U314 ( .A(n353), .B(n349), .CI(n351), .CO(n342), .S(n343) );
  CFA1X1 U315 ( .A(n374), .B(n355), .CI(n372), .CO(n344), .S(n345) );
  CFA1X1 U316 ( .A(n357), .B(n376), .CI(n378), .CO(n346), .S(n347) );
  CFA1X1 U317 ( .A(n741), .B(n380), .CI(n728), .CO(n348), .S(n349) );
  CFA1X1 U318 ( .A(n755), .B(n716), .CI(n695), .CO(n350), .S(n351) );
  CFA1X1 U320 ( .A(n705), .B(n660), .CI(n769), .CO(n354), .S(n355) );
  CHA1X1 U321 ( .A(n665), .B(n782), .CO(n356), .S(n357) );
  CFA1X1 U322 ( .A(n1014), .B(n1015), .CI(n1011), .CO(n358), .S(n359) );
  CFA1X1 U323 ( .A(n388), .B(n386), .CI(n365), .CO(n360), .S(n361) );
  CFA1X1 U324 ( .A(n390), .B(n367), .CI(n369), .CO(n362), .S(n363) );
  CFA1X1 U325 ( .A(n394), .B(n371), .CI(n392), .CO(n364), .S(n365) );
  CFA1X1 U326 ( .A(n373), .B(n375), .CI(n377), .CO(n366), .S(n367) );
  CFA1X1 U327 ( .A(n398), .B(n379), .CI(n396), .CO(n368), .S(n369) );
  CFA1X1 U328 ( .A(n402), .B(n400), .CI(n381), .CO(n370), .S(n371) );
  CFA1X1 U329 ( .A(n756), .B(n742), .CI(n729), .CO(n372), .S(n373) );
  CFA1X1 U330 ( .A(n770), .B(n717), .CI(n687), .CO(n374), .S(n375) );
  CFA1X1 U331 ( .A(n696), .B(n679), .CI(n672), .CO(n376), .S(n377) );
  CFA1X1 U332 ( .A(n706), .B(n783), .CI(n795), .CO(n378), .S(n379) );
  CHA1X1 U333 ( .A(a[13]), .B(n666), .CO(n380), .S(n381) );
  CFA1X1 U334 ( .A(n387), .B(n385), .CI(n406), .CO(n382), .S(n383) );
  CFA1X1 U335 ( .A(n391), .B(n389), .CI(n408), .CO(n384), .S(n385) );
  CFA1X1 U336 ( .A(n412), .B(n410), .CI(n393), .CO(n386), .S(n387) );
  CFA1X1 U337 ( .A(n397), .B(n395), .CI(n414), .CO(n388), .S(n389) );
  CFA1X1 U338 ( .A(n416), .B(n399), .CI(n401), .CO(n390), .S(n391) );
  CFA1X1 U339 ( .A(n422), .B(n420), .CI(n418), .CO(n392), .S(n393) );
  CFA1X1 U340 ( .A(n743), .B(n403), .CI(n424), .CO(n394), .S(n395) );
  CFA1X1 U341 ( .A(n757), .B(n697), .CI(n688), .CO(n396), .S(n397) );
  CFA1X1 U342 ( .A(n730), .B(n771), .CI(n784), .CO(n398), .S(n399) );
  CFA1X1 U343 ( .A(n718), .B(n680), .CI(n673), .CO(n400), .S(n401) );
  CHA1X1 U344 ( .A(n707), .B(n796), .CO(n402), .S(n403) );
  CFA1X1 U345 ( .A(n409), .B(n407), .CI(n428), .CO(n404), .S(n405) );
  CFA1X1 U346 ( .A(n413), .B(n430), .CI(n411), .CO(n406), .S(n407) );
  CFA1X1 U347 ( .A(n434), .B(n432), .CI(n415), .CO(n408), .S(n409) );
  CFA1X1 U348 ( .A(n423), .B(n436), .CI(n417), .CO(n410), .S(n411) );
  CFA1X1 U349 ( .A(n438), .B(n421), .CI(n419), .CO(n412), .S(n413) );
  CFA1X1 U350 ( .A(n425), .B(n440), .CI(n442), .CO(n414), .S(n415) );
  CFA1X1 U351 ( .A(n731), .B(n444), .CI(n719), .CO(n416), .S(n417) );
  CFA1X1 U352 ( .A(n758), .B(n689), .CI(n681), .CO(n418), .S(n419) );
  CFA1X1 U353 ( .A(n698), .B(n772), .CI(n797), .CO(n420), .S(n421) );
  CHA1X1 U355 ( .A(a[12]), .B(n708), .CO(n424), .S(n425) );
  CFA1X1 U356 ( .A(n431), .B(n429), .CI(n448), .CO(n426), .S(n427) );
  CFA1X1 U357 ( .A(n435), .B(n450), .CI(n433), .CO(n428), .S(n429) );
  CFA1X1 U358 ( .A(n454), .B(n452), .CI(n437), .CO(n430), .S(n431) );
  CFA1X1 U359 ( .A(n441), .B(n456), .CI(n443), .CO(n432), .S(n433) );
  CFA1X1 U360 ( .A(n460), .B(n439), .CI(n458), .CO(n434), .S(n435) );
  CFA1X1 U361 ( .A(n464), .B(n462), .CI(n445), .CO(n436), .S(n437) );
  CFA1X1 U362 ( .A(n773), .B(n759), .CI(n745), .CO(n438), .S(n439) );
  CFA1X1 U363 ( .A(n720), .B(n699), .CI(n690), .CO(n440), .S(n441) );
  CFA1X1 U364 ( .A(n732), .B(n786), .CI(n809), .CO(n442), .S(n443) );
  CHA1X1 U365 ( .A(n709), .B(n798), .CO(n444), .S(n445) );
  CFA1X1 U366 ( .A(n451), .B(n449), .CI(n468), .CO(n446), .S(n447) );
  CFA1X1 U367 ( .A(n455), .B(n470), .CI(n453), .CO(n448), .S(n449) );
  CFA1X1 U368 ( .A(n457), .B(n472), .CI(n474), .CO(n450), .S(n451) );
  CFA1X1 U369 ( .A(n459), .B(n461), .CI(n463), .CO(n452), .S(n453) );
  CFA1X1 U370 ( .A(n480), .B(n476), .CI(n478), .CO(n454), .S(n455) );
  CFA1X1 U371 ( .A(n746), .B(n465), .CI(n482), .CO(n456), .S(n457) );
  CFA1X1 U372 ( .A(n760), .B(n721), .CI(n700), .CO(n458), .S(n459) );
  CFA1X1 U373 ( .A(n733), .B(n787), .CI(n774), .CO(n460), .S(n461) );
  CFA1X1 U374 ( .A(n820), .B(n799), .CI(n810), .CO(n462), .S(n463) );
  CHA1X1 U375 ( .A(a[11]), .B(n710), .CO(n464), .S(n465) );
  CFA1X1 U376 ( .A(n471), .B(n469), .CI(n486), .CO(n466), .S(n467) );
  CFA1X1 U377 ( .A(n490), .B(n488), .CI(n473), .CO(n468), .S(n469) );
  CFA1X1 U378 ( .A(n477), .B(n475), .CI(n492), .CO(n470), .S(n471) );
  CFA1X1 U379 ( .A(n494), .B(n481), .CI(n479), .CO(n472), .S(n473) );
  CFA1X1 U380 ( .A(n483), .B(n496), .CI(n498), .CO(n474), .S(n475) );
  CFA1X1 U381 ( .A(n775), .B(n500), .CI(n747), .CO(n476), .S(n477) );
  CFA1X1 U382 ( .A(n734), .B(n811), .CI(n722), .CO(n478), .S(n479) );
  CFA1X1 U383 ( .A(n761), .B(n800), .CI(n788), .CO(n480), .S(n481) );
  CHA1X1 U384 ( .A(n711), .B(n821), .CO(n482), .S(n483) );
  CFA1X1 U385 ( .A(n489), .B(n487), .CI(n504), .CO(n484), .S(n485) );
  CFA1X1 U386 ( .A(n493), .B(n506), .CI(n491), .CO(n486), .S(n487) );
  CFA1X1 U387 ( .A(n499), .B(n508), .CI(n510), .CO(n488), .S(n489) );
  CFA1X1 U388 ( .A(n512), .B(n497), .CI(n495), .CO(n490), .S(n491) );
  CFA1X1 U389 ( .A(n516), .B(n514), .CI(n501), .CO(n492), .S(n493) );
  CFA1X1 U390 ( .A(n789), .B(n776), .CI(n748), .CO(n494), .S(n495) );
  CFA1X1 U391 ( .A(n762), .B(n822), .CI(n723), .CO(n496), .S(n497) );
  CFA1X1 U392 ( .A(n831), .B(n801), .CI(n812), .CO(n498), .S(n499) );
  CHA1X1 U393 ( .A(a[10]), .B(n735), .CO(n500), .S(n501) );
  CFA1X1 U394 ( .A(n507), .B(n505), .CI(n520), .CO(n502), .S(n503) );
  CFA1X1 U395 ( .A(n511), .B(n509), .CI(n522), .CO(n504), .S(n505) );
  CFA1X1 U396 ( .A(n513), .B(n524), .CI(n515), .CO(n506), .S(n507) );
  CFA1X1 U397 ( .A(n530), .B(n526), .CI(n528), .CO(n508), .S(n509) );
  CFA1X1 U398 ( .A(n832), .B(n517), .CI(n532), .CO(n510), .S(n511) );
  CFA1X1 U399 ( .A(n749), .B(n802), .CI(n986), .CO(n512), .S(n513) );
  CFA1X1 U400 ( .A(n777), .B(n823), .CI(n813), .CO(n514), .S(n515) );
  CHA1X1 U401 ( .A(n736), .B(n790), .CO(n516), .S(n517) );
  CFA1X1 U402 ( .A(n523), .B(n521), .CI(n536), .CO(n518), .S(n519) );
  CFA1X1 U403 ( .A(n540), .B(n538), .CI(n525), .CO(n520), .S(n521) );
  CFA1X1 U404 ( .A(n529), .B(n527), .CI(n531), .CO(n522), .S(n523) );
  CFA1X1 U405 ( .A(n533), .B(n542), .CI(n544), .CO(n524), .S(n525) );
  CFA1X1 U406 ( .A(n833), .B(n546), .CI(n764), .CO(n526), .S(n527) );
  CFA1X1 U407 ( .A(n778), .B(n791), .CI(n824), .CO(n528), .S(n529) );
  CFA1X1 U408 ( .A(n814), .B(n841), .CI(n803), .CO(n530), .S(n531) );
  CFA1X1 U410 ( .A(n539), .B(n537), .CI(n550), .CO(n534), .S(n535) );
  CFA1X1 U411 ( .A(n554), .B(n552), .CI(n541), .CO(n536), .S(n537) );
  CFA1X1 U412 ( .A(n556), .B(n545), .CI(n543), .CO(n538), .S(n539) );
  CFA1X1 U413 ( .A(n560), .B(n558), .CI(n547), .CO(n540), .S(n541) );
  CFA1X1 U414 ( .A(n825), .B(n804), .CI(n765), .CO(n542), .S(n543) );
  CFA1X1 U415 ( .A(n834), .B(n792), .CI(n842), .CO(n544), .S(n545) );
  CHA1X1 U416 ( .A(n779), .B(n815), .CO(n546), .S(n547) );
  CFA1X1 U417 ( .A(n553), .B(n551), .CI(n564), .CO(n548), .S(n549) );
  CFA1X1 U418 ( .A(n557), .B(n566), .CI(n555), .CO(n550), .S(n551) );
  CFA1X1 U419 ( .A(n570), .B(n559), .CI(n568), .CO(n552), .S(n553) );
  CFA1X1 U420 ( .A(n843), .B(n561), .CI(n572), .CO(n554), .S(n555) );
  CFA1X1 U421 ( .A(n816), .B(n826), .CI(n850), .CO(n556), .S(n557) );
  CFA1X1 U422 ( .A(n835), .B(n805), .CI(n793), .CO(n558), .S(n559) );
  CHA1X1 U423 ( .A(a[8]), .B(n780), .CO(n560), .S(n561) );
  CFA1X1 U424 ( .A(n567), .B(n565), .CI(n576), .CO(n562), .S(n563) );
  CFA1X1 U425 ( .A(n571), .B(n578), .CI(n569), .CO(n564), .S(n565) );
  CFA1X1 U426 ( .A(n573), .B(n580), .CI(n582), .CO(n566), .S(n567) );
  CFA1X1 U427 ( .A(n817), .B(n584), .CI(n806), .CO(n568), .S(n569) );
  CFA1X1 U428 ( .A(n836), .B(n827), .CI(n851), .CO(n570), .S(n571) );
  CHA1X1 U429 ( .A(n844), .B(n794), .CO(n572), .S(n573) );
  CFA1X1 U430 ( .A(n579), .B(n577), .CI(n588), .CO(n574), .S(n575) );
  CFA1X1 U431 ( .A(n583), .B(n590), .CI(n581), .CO(n576), .S(n577) );
  CFA1X1 U432 ( .A(n594), .B(n592), .CI(n585), .CO(n578), .S(n579) );
  CFA1X1 U433 ( .A(n845), .B(n828), .CI(n818), .CO(n580), .S(n581) );
  CFA1X1 U434 ( .A(n837), .B(n858), .CI(n807), .CO(n582), .S(n583) );
  CHA1X1 U435 ( .A(a[7]), .B(n852), .CO(n584), .S(n585) );
  CFA1X1 U436 ( .A(n591), .B(n589), .CI(n598), .CO(n586), .S(n587) );
  CFA1X1 U437 ( .A(n602), .B(n593), .CI(n600), .CO(n588), .S(n589) );
  CFA1X1 U438 ( .A(n846), .B(n595), .CI(n604), .CO(n590), .S(n591) );
  CFA1X1 U439 ( .A(n859), .B(n829), .CI(n853), .CO(n592), .S(n593) );
  CHA1X1 U440 ( .A(n838), .B(n819), .CO(n594), .S(n595) );
  CFA1X1 U441 ( .A(n601), .B(n599), .CI(n608), .CO(n596), .S(n597) );
  CFA1X1 U442 ( .A(n605), .B(n603), .CI(n610), .CO(n598), .S(n599) );
  CFA1X1 U443 ( .A(n854), .B(n612), .CI(n847), .CO(n600), .S(n601) );
  CFA1X1 U444 ( .A(n865), .B(n860), .CI(n830), .CO(n602), .S(n603) );
  CHA1X1 U445 ( .A(a[6]), .B(n839), .CO(n604), .S(n605) );
  CFA1X1 U446 ( .A(n611), .B(n609), .CI(n616), .CO(n606), .S(n607) );
  CFA1X1 U447 ( .A(n620), .B(n618), .CI(n613), .CO(n608), .S(n609) );
  CFA1X1 U448 ( .A(n855), .B(n866), .CI(n861), .CO(n610), .S(n611) );
  CHA1X1 U449 ( .A(n840), .B(n848), .CO(n612), .S(n613) );
  CFA1X1 U450 ( .A(n624), .B(n617), .CI(n619), .CO(n614), .S(n615) );
  CFA1X1 U451 ( .A(n862), .B(n621), .CI(n626), .CO(n616), .S(n617) );
  CFA1X1 U452 ( .A(n867), .B(n856), .CI(n849), .CO(n618), .S(n619) );
  CHA1X1 U453 ( .A(a[5]), .B(n871), .CO(n620), .S(n621) );
  CFA1X1 U454 ( .A(n627), .B(n625), .CI(n630), .CO(n622), .S(n623) );
  CFA1X1 U455 ( .A(n868), .B(n632), .CI(n863), .CO(n624), .S(n625) );
  CHA1X1 U456 ( .A(n872), .B(n857), .CO(n626), .S(n627) );
  CFA1X1 U457 ( .A(n636), .B(n631), .CI(n633), .CO(n628), .S(n629) );
  CFA1X1 U458 ( .A(n876), .B(n869), .CI(n864), .CO(n630), .S(n631) );
  CHA1X1 U459 ( .A(a[4]), .B(n873), .CO(n632), .S(n633) );
  CFA1X1 U460 ( .A(n877), .B(n637), .CI(n640), .CO(n634), .S(n635) );
  CHA1X1 U461 ( .A(n874), .B(n870), .CO(n636), .S(n637) );
  CFA1X1 U462 ( .A(n880), .B(n642), .CI(n878), .CO(n638), .S(n639) );
  CHA1X1 U463 ( .A(a[3]), .B(n875), .CO(n640), .S(n641) );
  CHA1X1 U464 ( .A(n881), .B(n879), .CO(n642), .S(n643) );
  CFD1QXL clk_r_REG49_S1 ( .D(n997), .CP(n1058), .Q(n1053) );
  CFD1QXL clk_r_REG48_S1 ( .D(n177), .CP(n1058), .Q(n1052) );
  CFD1QXL clk_r_REG0_S1 ( .D(n257), .CP(n1058), .Q(n1027) );
  CFD1QXL clk_r_REG44_S1 ( .D(n165), .CP(n1058), .Q(n1034) );
  CFD1QXL clk_r_REG43_S1 ( .D(n166), .CP(n1058), .Q(n1033) );
  CFD1QXL clk_r_REG6_S1 ( .D(n259), .CP(n1058), .Q(n1026) );
  CFD1QXL clk_r_REG36_S1 ( .D(n73), .CP(n1058), .Q(n1035) );
  CFD1QXL clk_r_REG41_S1 ( .D(n75), .CP(n1058), .Q(n1032) );
  CFD1QXL clk_r_REG47_S1 ( .D(n76), .CP(n1058), .Q(n1031) );
  CFD1QXL clk_r_REG1_S1 ( .D(n240), .CP(n1058), .Q(n1028) );
  CFD1QXL clk_r_REG46_S1 ( .D(n180), .CP(n1058), .Q(n1051) );
  CFD1QXL clk_r_REG38_S1 ( .D(n160), .CP(n1058), .Q(n1036) );
  CFD1QXL clk_r_REG37_S1 ( .D(n161), .CP(n1058), .Q(n1030) );
  CFD1QXL clk_r_REG27_S1 ( .D(n118), .CP(n1058), .Q(n1046) );
  CFD1QXL clk_r_REG4_S1 ( .D(n285), .CP(n1058), .Q(n1024) );
  CFD1QXL clk_r_REG35_S1 ( .D(n139), .CP(n1058), .Q(n1040) );
  CFD1QXL clk_r_REG21_S1 ( .D(n108), .CP(n1058), .Q(n1049) );
  CFD1QXL clk_r_REG11_S1 ( .D(n310), .CP(n1058), .Q(n1022) );
  CFD1QXL clk_r_REG9_S1 ( .D(n336), .CP(n1058), .Q(n1019) );
  CFD1QXL clk_r_REG7_S1 ( .D(n360), .CP(n1058), .Q(n1016) );
  CFD1QXL clk_r_REG16_S1 ( .D(n384), .CP(n1058), .Q(n1011) );
  CFD1QXL clk_r_REG5_S1 ( .D(n287), .CP(n1058), .Q(n1023) );
  CFD1QXL clk_r_REG2_S1 ( .D(n313), .CP(n1058), .Q(n1020) );
  CFD1QXL clk_r_REG13_S1 ( .D(n339), .CP(n1058), .Q(n1017) );
  CFD1QXL clk_r_REG58_S1 ( .D(n363), .CP(n1058), .Q(n1014) );
  CFD1QXL clk_r_REG26_S1 ( .D(n119), .CP(n1058), .Q(n1045) );
  CFD1QXL clk_r_REG24_S1 ( .D(n124), .CP(n1058), .Q(n1044) );
  CFD1QXL clk_r_REG32_S1 ( .D(n152), .CP(n1058), .Q(n1038) );
  CFD1QXL clk_r_REG28_S1 ( .D(n137), .CP(n1058), .Q(n1041) );
  CFD1QXL clk_r_REG39_S1 ( .D(n157), .CP(n1058), .Q(n1037) );
  CFD1QXL clk_r_REG18_S1 ( .D(n383), .CP(n1058), .Q(n1012) );
  CFD1QXL clk_r_REG15_S1 ( .D(n405), .CP(n1058), .Q(n1009) );
  CFD1QXL clk_r_REG19_S1 ( .D(n111), .CP(n1058), .Q(n1047) );
  CFD1QXL clk_r_REG17_S1 ( .D(n382), .CP(n1058), .Q(n1013) );
  CFD1QXL clk_r_REG14_S1 ( .D(n404), .CP(n1058), .Q(n1010) );
  CFD1QXL clk_r_REG22_S1 ( .D(n107), .CP(n1058), .Q(n1050) );
  CFD1QXL clk_r_REG33_S1 ( .D(n994), .CP(n1058), .Q(n1055) );
  CFD1QXL clk_r_REG29_S1 ( .D(n995), .CP(n1058), .Q(n1056) );
  CFD1QXL clk_r_REG20_S1 ( .D(n110), .CP(n1058), .Q(n1048) );
  CFD1QXL clk_r_REG34_S1 ( .D(n140), .CP(n1058), .Q(n1039) );
  CFD1QXL clk_r_REG25_S1 ( .D(n996), .CP(n1058), .Q(n1057) );
  CFD1QXL clk_r_REG40_S1 ( .D(n1000), .CP(n1058), .Q(n1054) );
  CFD1QXL clk_r_REG23_S1 ( .D(n426), .CP(n1058), .Q(n1008) );
  CFD1QXL clk_r_REG8_S1 ( .D(n361), .CP(n1058), .Q(n1015) );
  CFD1QXL clk_r_REG3_S1 ( .D(n284), .CP(n1058), .Q(n1025) );
  CFD1QXL clk_r_REG12_S1 ( .D(n311), .CP(n1058), .Q(n1021) );
  CFD1QXL clk_r_REG30_S1 ( .D(n130), .CP(n1058), .Q(n1042) );
  CFD1QXL clk_r_REG31_S1 ( .D(n129), .CP(n1058), .Q(n1043) );
  CFD1QXL clk_r_REG10_S1 ( .D(n337), .CP(n1058), .Q(n1018) );
  CFD1QX2 clk_r_REG42_S1 ( .D(n168), .CP(n1058), .Q(n1029) );
  CNR2XL U754 ( .A(n32), .B(n48), .Z(n857) );
  CNR2XL U755 ( .A(n32), .B(n38), .Z(n882) );
  CNR2XL U756 ( .A(n32), .B(n50), .Z(n849) );
  CNR2XL U757 ( .A(n32), .B(n912), .Z(n819) );
  CNR2XL U758 ( .A(n32), .B(n911), .Z(n807) );
  CNR2X1 U759 ( .A(n32), .B(n22), .Z(n690) );
  COND1X1 U760 ( .A(n1043), .B(n133), .C(n1042), .Z(n128) );
  CIVXL U761 ( .A(n126), .Z(n125) );
  CNIVX1 U762 ( .A(n763), .Z(n986) );
  CNIVX1 U763 ( .A(n738), .Z(n987) );
  CNR2X1 U764 ( .A(n40), .B(n22), .Z(n686) );
  CIVX1 U765 ( .A(b[22]), .Z(n22) );
  CFA1X1 U766 ( .A(n686), .B(n678), .CI(n671), .CO(n352), .S(n353) );
  CNR2X1 U767 ( .A(n36), .B(n24), .Z(n671) );
  CNR2X1 U768 ( .A(n36), .B(n26), .Z(n658) );
  CNR2X1 U769 ( .A(n32), .B(n20), .Z(n711) );
  CIVX3 U770 ( .A(b[17]), .Z(n17) );
  CFA1XL U771 ( .A(n744), .B(n785), .CI(n808), .CO(n422), .S(n423) );
  CHA1X1 U772 ( .A(a[9]), .B(n750), .CO(n532), .S(n533) );
  CNR2X1 U773 ( .A(n32), .B(n17), .Z(n750) );
  CNR2IXL U774 ( .B(b[11]), .A(n17), .Z(n739) );
  CIVX3 U775 ( .A(b[11]), .Z(n54) );
  CNIVX1 U776 ( .A(n989), .Z(product[12]) );
  CNIVX1 U777 ( .A(n1090), .Z(n989) );
  CNIVX1 U778 ( .A(n991), .Z(product[14]) );
  CNIVX1 U779 ( .A(n1089), .Z(n991) );
  CNIVX1 U780 ( .A(n1091), .Z(product[11]) );
  CIVX4 U781 ( .A(b[2]), .Z(n36) );
  CHA1XL U782 ( .A(a[2]), .B(n883), .CO(n644), .S(n645) );
  CFA1XL U783 ( .A(n726), .B(n669), .CI(n658), .CO(n300), .S(n301) );
  CIVX1 U784 ( .A(n1038), .Z(n150) );
  COND1X2 U785 ( .A(n102), .B(n104), .C(n103), .Z(n101) );
  CANR1X2 U786 ( .A(n105), .B(n113), .C(n106), .Z(n104) );
  COND1X2 U787 ( .A(n94), .B(n96), .C(n95), .Z(n93) );
  CANR1X2 U788 ( .A(n1007), .B(n101), .C(n98), .Z(n96) );
  CNR2XL U789 ( .A(n36), .B(n46), .Z(n862) );
  CNR2XL U790 ( .A(n36), .B(n50), .Z(n847) );
  CNR2XL U791 ( .A(n36), .B(n40), .Z(n877) );
  COR2XL U792 ( .A(n32), .B(n36), .Z(n1002) );
  CNR2XL U793 ( .A(n36), .B(n52), .Z(n838) );
  CNR2XL U794 ( .A(n36), .B(n48), .Z(n855) );
  CNR2XL U795 ( .A(n36), .B(n28), .Z(n649) );
  CNR2XL U796 ( .A(n36), .B(n911), .Z(n805) );
  CNR2XL U797 ( .A(n36), .B(n27), .Z(n653) );
  CNR2XL U798 ( .A(n34), .B(n36), .Z(n883) );
  CNR2XL U799 ( .A(n36), .B(n15), .Z(n778) );
  CNR2XL U800 ( .A(n36), .B(n16), .Z(n763) );
  CANR1X2 U801 ( .A(n202), .B(n1006), .C(n199), .Z(n197) );
  COND1X1 U802 ( .A(n203), .B(n205), .C(n204), .Z(n202) );
  CIVXL U803 ( .A(n181), .Z(n180) );
  CANR1X1 U804 ( .A(n999), .B(n186), .C(n183), .Z(n181) );
  COND1X1 U805 ( .A(n147), .B(n159), .C(n148), .Z(n146) );
  CANR1X1 U806 ( .A(n1036), .B(n1029), .C(n1030), .Z(n159) );
  COND1X2 U807 ( .A(n114), .B(n126), .C(n115), .Z(n113) );
  CANR1X2 U808 ( .A(n146), .B(n127), .C(n128), .Z(n126) );
  CNR2XL U809 ( .A(n38), .B(n27), .Z(n652) );
  CNR2XL U810 ( .A(n50), .B(n19), .Z(n714) );
  CNR2XL U811 ( .A(n36), .B(n25), .Z(n664) );
  CNR2XL U812 ( .A(n52), .B(n18), .Z(n726) );
  CNR2XL U813 ( .A(n42), .B(n25), .Z(n661) );
  CNR2X1 U814 ( .A(n38), .B(n40), .Z(n876) );
  CNR2XL U815 ( .A(n912), .B(n17), .Z(n738) );
  CNR2XL U816 ( .A(n34), .B(n28), .Z(n650) );
  CNR2XL U817 ( .A(n46), .B(n910), .Z(n787) );
  CND2XL U818 ( .A(n1056), .B(n225), .Z(n132) );
  CEOXL U819 ( .A(n197), .B(n80), .Z(product[7]) );
  CANR1XL U820 ( .A(n210), .B(n1003), .C(n207), .Z(n205) );
  CNR2XL U821 ( .A(n38), .B(n912), .Z(n816) );
  CNR2X1 U822 ( .A(n32), .B(n27), .Z(n655) );
  CNR2XL U823 ( .A(n42), .B(n15), .Z(n775) );
  CNR2XL U824 ( .A(n40), .B(n52), .Z(n836) );
  CNR2XL U825 ( .A(n50), .B(n42), .Z(n844) );
  CNR2XL U826 ( .A(n36), .B(n912), .Z(n817) );
  CNR2X1 U827 ( .A(n34), .B(n23), .Z(n680) );
  CNR2XL U828 ( .A(n32), .B(n52), .Z(n840) );
  CNR2XL U829 ( .A(n46), .B(n42), .Z(n859) );
  CNR2XL U830 ( .A(n38), .B(n44), .Z(n867) );
  CNR2XL U831 ( .A(n32), .B(n40), .Z(n879) );
  CNR2XL U832 ( .A(n40), .B(n912), .Z(n815) );
  CNR2XL U833 ( .A(n36), .B(n44), .Z(n868) );
  CNR2XL U834 ( .A(n911), .B(n52), .Z(n797) );
  CNR2XL U835 ( .A(n46), .B(n52), .Z(n833) );
  CNR2XL U836 ( .A(n44), .B(n42), .Z(n865) );
  CNR2XL U837 ( .A(n42), .B(n52), .Z(n835) );
  CNR2XL U838 ( .A(n32), .B(n44), .Z(n870) );
  CNR2XL U839 ( .A(n32), .B(n30), .Z(n646) );
  CNR2XL U840 ( .A(n36), .B(n38), .Z(n880) );
  CIVX2 U841 ( .A(b[13]), .Z(n911) );
  CIVX2 U842 ( .A(b[15]), .Z(n15) );
  CIVX3 U843 ( .A(b[9]), .Z(n50) );
  CND2XL U844 ( .A(n885), .B(a[1]), .Z(n213) );
  CND2XL U845 ( .A(n999), .B(n185), .Z(n77) );
  CNR2XL U846 ( .A(n427), .B(n446), .Z(n107) );
  CNR2XL U847 ( .A(n447), .B(n466), .Z(n110) );
  CNR2XL U848 ( .A(n467), .B(n484), .Z(n118) );
  CNR2XL U849 ( .A(n162), .B(n165), .Z(n160) );
  CNR2XL U850 ( .A(n503), .B(n518), .Z(n129) );
  CNR2XL U851 ( .A(n535), .B(n548), .Z(n139) );
  CND2XL U852 ( .A(n485), .B(n502), .Z(n124) );
  CND2XL U853 ( .A(n503), .B(n518), .Z(n130) );
  CND2XL U854 ( .A(n998), .B(n174), .Z(n75) );
  CND2XL U855 ( .A(n535), .B(n548), .Z(n140) );
  CND2XL U856 ( .A(n549), .B(n562), .Z(n152) );
  CND2XL U857 ( .A(n997), .B(n179), .Z(n76) );
  CND2XL U858 ( .A(n519), .B(n534), .Z(n137) );
  CND2IXL U859 ( .B(n162), .A(n163), .Z(n73) );
  CIVXL U860 ( .A(n179), .Z(n177) );
  CND2XL U861 ( .A(n233), .B(n188), .Z(n78) );
  CND2XL U862 ( .A(n235), .B(n196), .Z(n80) );
  CND2XL U863 ( .A(n1001), .B(n193), .Z(n79) );
  CND2XL U864 ( .A(n575), .B(n586), .Z(n163) );
  CND2XL U865 ( .A(n563), .B(n574), .Z(n157) );
  CND2XL U866 ( .A(n237), .B(n204), .Z(n82) );
  CND2XL U867 ( .A(n1003), .B(n209), .Z(n83) );
  CND2XL U868 ( .A(n1006), .B(n201), .Z(n81) );
  CNR2XL U869 ( .A(n48), .B(n54), .Z(n822) );
  CNR2XL U870 ( .A(n34), .B(n44), .Z(n869) );
  CNR2XL U871 ( .A(n46), .B(n54), .Z(n823) );
  CNR2XL U872 ( .A(n36), .B(n910), .Z(n792) );
  CNR2XL U873 ( .A(n40), .B(n54), .Z(n826) );
  CNR2XL U874 ( .A(n34), .B(n48), .Z(n856) );
  CNR2XL U875 ( .A(n34), .B(n24), .Z(n672) );
  CNR2XL U876 ( .A(n36), .B(n23), .Z(n679) );
  CNR2XL U877 ( .A(n40), .B(n21), .Z(n696) );
  CNR2XL U878 ( .A(n52), .B(n17), .Z(n740) );
  CNR2XL U879 ( .A(n34), .B(n26), .Z(n659) );
  CNR2XL U880 ( .A(n46), .B(n18), .Z(n729) );
  CNR2XL U881 ( .A(n48), .B(n17), .Z(n742) );
  CNR2XL U882 ( .A(n50), .B(n16), .Z(n756) );
  CNR2XL U883 ( .A(n46), .B(n23), .Z(n674) );
  CNR2XL U884 ( .A(n50), .B(n21), .Z(n691) );
  CNR2XL U885 ( .A(n40), .B(n26), .Z(n656) );
  CNR2XL U886 ( .A(n54), .B(n19), .Z(n712) );
  CNR2XL U887 ( .A(n50), .B(n54), .Z(n821) );
  CNR2XL U888 ( .A(n34), .B(n15), .Z(n779) );
  CNR2XL U889 ( .A(n54), .B(n16), .Z(n754) );
  CNR2XL U890 ( .A(n42), .B(n22), .Z(n685) );
  CNR2XL U891 ( .A(n46), .B(n21), .Z(n693) );
  CNR2XL U892 ( .A(n38), .B(n22), .Z(n687) );
  CNR2XL U893 ( .A(n44), .B(n19), .Z(n717) );
  CEOXL U894 ( .A(n213), .B(n1002), .Z(product[3]) );
  CNR2XL U895 ( .A(n38), .B(n17), .Z(n747) );
  CNR2XL U896 ( .A(n40), .B(n17), .Z(n746) );
  CNR2XL U897 ( .A(n38), .B(n910), .Z(n791) );
  CNR2XL U898 ( .A(n44), .B(n54), .Z(n824) );
  CNR2XL U899 ( .A(n38), .B(n54), .Z(n827) );
  CNR2XL U900 ( .A(n48), .B(n21), .Z(n692) );
  CNR2XL U901 ( .A(n52), .B(n19), .Z(n713) );
  CNR2XL U902 ( .A(n911), .B(n910), .Z(n781) );
  CNR2XL U903 ( .A(n44), .B(n17), .Z(n744) );
  CNR2XL U904 ( .A(n50), .B(n910), .Z(n785) );
  CNR2XL U905 ( .A(n54), .B(n912), .Z(n808) );
  CNR2XL U906 ( .A(n36), .B(n22), .Z(n688) );
  CNR2XL U907 ( .A(n38), .B(n21), .Z(n697) );
  CNR2XL U908 ( .A(n48), .B(n16), .Z(n757) );
  CNR2XL U909 ( .A(n42), .B(n20), .Z(n706) );
  CNR2XL U910 ( .A(n54), .B(n910), .Z(n783) );
  CNR2XL U911 ( .A(n46), .B(n19), .Z(n716) );
  CNR2XL U912 ( .A(n44), .B(n21), .Z(n694) );
  CNR2XL U913 ( .A(n50), .B(n18), .Z(n727) );
  CNR2XL U914 ( .A(n34), .B(n25), .Z(n665) );
  CNR2XL U915 ( .A(n912), .B(n910), .Z(n782) );
  CNR2XL U916 ( .A(n32), .B(n910), .Z(n794) );
  CNR2XL U917 ( .A(n34), .B(n911), .Z(n806) );
  CNR2XL U918 ( .A(n38), .B(n26), .Z(n657) );
  CNR2XL U919 ( .A(n46), .B(n22), .Z(n683) );
  CNR2XL U920 ( .A(n54), .B(n18), .Z(n725) );
  CNR2XL U921 ( .A(n42), .B(n19), .Z(n718) );
  CNR2XL U922 ( .A(n42), .B(n18), .Z(n731) );
  CNR2XL U923 ( .A(n40), .B(n19), .Z(n719) );
  CNR2XL U924 ( .A(n34), .B(n912), .Z(n818) );
  CNR2XL U925 ( .A(n36), .B(n54), .Z(n828) );
  CNR2XL U926 ( .A(n34), .B(n22), .Z(n689) );
  CNR2XL U927 ( .A(n46), .B(n16), .Z(n758) );
  CNR2XL U928 ( .A(n34), .B(n50), .Z(n848) );
  CNR2XL U929 ( .A(n911), .B(n17), .Z(n737) );
  CNR2XL U930 ( .A(n44), .B(n24), .Z(n667) );
  CNR2XL U931 ( .A(n52), .B(n20), .Z(n701) );
  CNR2XL U932 ( .A(n32), .B(n34), .Z(n885) );
  CNR2XL U933 ( .A(n48), .B(n19), .Z(n715) );
  CNR2XL U934 ( .A(n34), .B(n54), .Z(n829) );
  CNR2XL U935 ( .A(n34), .B(n38), .Z(n881) );
  CNR2XL U936 ( .A(n36), .B(n20), .Z(n709) );
  CNR2XL U937 ( .A(n38), .B(n25), .Z(n663) );
  CNR2XL U938 ( .A(n34), .B(n46), .Z(n863) );
  CNR2XL U939 ( .A(n34), .B(n16), .Z(n764) );
  CNR2XL U940 ( .A(n46), .B(n17), .Z(n743) );
  CNR2XL U941 ( .A(n910), .B(n15), .Z(n766) );
  CNR2XL U942 ( .A(n32), .B(n54), .Z(n830) );
  CNR2XL U943 ( .A(n50), .B(n17), .Z(n741) );
  CNR2XL U944 ( .A(n48), .B(n18), .Z(n728) );
  CNR2XL U945 ( .A(n34), .B(n910), .Z(n793) );
  CNR2XL U946 ( .A(n36), .B(n21), .Z(n698) );
  CNR2XL U947 ( .A(n44), .B(n18), .Z(n730) );
  CNR2XL U948 ( .A(n910), .B(n52), .Z(n784) );
  CNR2XL U949 ( .A(n34), .B(n42), .Z(n874) );
  CNR2XL U950 ( .A(n32), .B(n18), .Z(n736) );
  CNR2XL U951 ( .A(n40), .B(n910), .Z(n790) );
  CNR2XL U952 ( .A(n34), .B(n29), .Z(n647) );
  CNR2XL U953 ( .A(n912), .B(n18), .Z(n724) );
  CEO3X1 U954 ( .A(n724), .B(n280), .C(n278), .Z(n248) );
  CNR2XL U955 ( .A(n911), .B(n16), .Z(n752) );
  CNR2XL U956 ( .A(n910), .B(n16), .Z(n751) );
  CEO3X1 U957 ( .A(n661), .B(n652), .C(n656), .Z(n251) );
  CNR2XL U958 ( .A(n48), .B(n22), .Z(n682) );
  CEO3X1 U959 ( .A(n737), .B(n691), .C(n712), .Z(n249) );
  CNR2XL U960 ( .A(n34), .B(n40), .Z(n878) );
  CIVX4 U961 ( .A(b[3]), .Z(n38) );
  CIVX4 U962 ( .A(b[4]), .Z(n40) );
  CNR2XL U963 ( .A(n132), .B(n1043), .Z(n127) );
  CIVX4 U964 ( .A(b[6]), .Z(n44) );
  CIVX4 U965 ( .A(b[5]), .Z(n42) );
  CIVX4 U966 ( .A(b[7]), .Z(n46) );
  CIVX4 U967 ( .A(b[8]), .Z(n48) );
  CIVX4 U968 ( .A(b[10]), .Z(n52) );
  CIVX4 U969 ( .A(\b[0] ), .Z(n32) );
  CIVX3 U970 ( .A(b[12]), .Z(n912) );
  CENX1 U971 ( .A(n993), .B(n85), .Z(product[31]) );
  CENX1 U972 ( .A(n1028), .B(n254), .Z(n993) );
  CND2XL U973 ( .A(n220), .B(n1047), .Z(n65) );
  CNR2XL U974 ( .A(n40), .B(n42), .Z(n871) );
  CIVX1 U975 ( .A(b[28]), .Z(n28) );
  CIVXL U976 ( .A(n1041), .Z(n135) );
  CND2IXL U977 ( .B(n212), .A(n213), .Z(n84) );
  CENX1 U978 ( .A(n77), .B(n186), .Z(product[10]) );
  COND1XL U979 ( .A(n181), .B(n169), .C(n170), .Z(n168) );
  CND2X1 U980 ( .A(n998), .B(n997), .Z(n169) );
  CANR1XL U981 ( .A(n177), .B(n998), .C(n172), .Z(n170) );
  COND1XL U982 ( .A(n166), .B(n162), .C(n163), .Z(n161) );
  COR2X1 U983 ( .A(n549), .B(n562), .Z(n994) );
  CND2XL U984 ( .A(n427), .B(n446), .Z(n108) );
  CND2XL U985 ( .A(n467), .B(n484), .Z(n119) );
  CND2XL U986 ( .A(n447), .B(n466), .Z(n111) );
  COR2X1 U987 ( .A(n519), .B(n534), .Z(n995) );
  COR2X1 U988 ( .A(n485), .B(n502), .Z(n996) );
  CANR1XL U989 ( .A(n194), .B(n1001), .C(n191), .Z(n189) );
  COND1XL U990 ( .A(n195), .B(n197), .C(n196), .Z(n194) );
  COND1XL U991 ( .A(n187), .B(n189), .C(n188), .Z(n186) );
  CNR2X1 U992 ( .A(n575), .B(n586), .Z(n162) );
  CENX1 U993 ( .A(n79), .B(n194), .Z(product[8]) );
  CNR2X1 U994 ( .A(n587), .B(n596), .Z(n165) );
  CEOXL U995 ( .A(n189), .B(n78), .Z(product[9]) );
  COR2X1 U996 ( .A(n607), .B(n614), .Z(n997) );
  COR2X1 U997 ( .A(n597), .B(n606), .Z(n998) );
  CND2X1 U998 ( .A(n597), .B(n606), .Z(n174) );
  CND2X1 U999 ( .A(n615), .B(n622), .Z(n185) );
  CND2X1 U1000 ( .A(n607), .B(n614), .Z(n179) );
  COR2X1 U1001 ( .A(n615), .B(n622), .Z(n999) );
  CND2X1 U1002 ( .A(n587), .B(n596), .Z(n166) );
  COR2X1 U1003 ( .A(n563), .B(n574), .Z(n1000) );
  CENX1 U1004 ( .A(n81), .B(n202), .Z(product[6]) );
  CENX1 U1005 ( .A(n93), .B(n60), .Z(product[27]) );
  CND2X1 U1006 ( .A(n1005), .B(n92), .Z(n60) );
  CNR2X1 U1007 ( .A(n635), .B(n638), .Z(n195) );
  CNR2X1 U1008 ( .A(n623), .B(n628), .Z(n187) );
  CEOXL U1009 ( .A(n205), .B(n82), .Z(product[5]) );
  CND2X1 U1010 ( .A(n629), .B(n634), .Z(n193) );
  CND2X1 U1011 ( .A(n635), .B(n638), .Z(n196) );
  CND2X1 U1012 ( .A(n623), .B(n628), .Z(n188) );
  COR2X1 U1013 ( .A(n629), .B(n634), .Z(n1001) );
  CENX1 U1014 ( .A(n83), .B(n210), .Z(product[4]) );
  CNR2X1 U1015 ( .A(n213), .B(n1002), .Z(n210) );
  CNR2X1 U1016 ( .A(n40), .B(n46), .Z(n860) );
  CNR2X1 U1017 ( .A(n42), .B(n24), .Z(n668) );
  CNR2X1 U1018 ( .A(n40), .B(n48), .Z(n853) );
  CNR2X1 U1019 ( .A(n48), .B(n911), .Z(n799) );
  CNR2X1 U1020 ( .A(n50), .B(n912), .Z(n810) );
  CNR2X1 U1021 ( .A(n54), .B(n52), .Z(n820) );
  CNR2X1 U1022 ( .A(n38), .B(n911), .Z(n804) );
  CNR2X1 U1023 ( .A(n32), .B(n16), .Z(n765) );
  CNR2X1 U1024 ( .A(n54), .B(n42), .Z(n825) );
  CNR2X1 U1025 ( .A(n912), .B(n15), .Z(n768) );
  CNR2X1 U1026 ( .A(n40), .B(n23), .Z(n677) );
  CENX1 U1027 ( .A(n101), .B(n62), .Z(product[25]) );
  CND2X1 U1028 ( .A(n1007), .B(n100), .Z(n62) );
  CNR2X1 U1029 ( .A(n911), .B(n42), .Z(n802) );
  CNR2X1 U1030 ( .A(n34), .B(n17), .Z(n749) );
  CNR2X1 U1031 ( .A(n48), .B(n50), .Z(n841) );
  CNR2X1 U1032 ( .A(n40), .B(n911), .Z(n803) );
  CNR2X1 U1033 ( .A(n912), .B(n42), .Z(n814) );
  CNR2X1 U1034 ( .A(n44), .B(n15), .Z(n774) );
  CNR2X1 U1035 ( .A(n38), .B(n18), .Z(n733) );
  CNR2X1 U1036 ( .A(n42), .B(n23), .Z(n676) );
  CNR2X1 U1037 ( .A(n46), .B(n48), .Z(n850) );
  CNR2X1 U1038 ( .A(n52), .B(n15), .Z(n770) );
  CNR2X1 U1039 ( .A(n44), .B(n48), .Z(n851) );
  CNR2X1 U1040 ( .A(n643), .B(n644), .Z(n203) );
  CNR2X1 U1041 ( .A(n36), .B(n19), .Z(n721) );
  CNR2X1 U1042 ( .A(n42), .B(n16), .Z(n760) );
  CNR2X1 U1043 ( .A(n32), .B(n21), .Z(n700) );
  CNR2X1 U1044 ( .A(n48), .B(n52), .Z(n832) );
  CNR2X1 U1045 ( .A(n44), .B(n911), .Z(n801) );
  CNR2X1 U1046 ( .A(n46), .B(n912), .Z(n812) );
  CNR2X1 U1047 ( .A(n50), .B(n52), .Z(n831) );
  CNR2X1 U1048 ( .A(n46), .B(n50), .Z(n842) );
  CNR2X1 U1049 ( .A(n44), .B(n52), .Z(n834) );
  CNR2X1 U1050 ( .A(n40), .B(n24), .Z(n669) );
  CNR2X1 U1051 ( .A(n44), .B(n46), .Z(n858) );
  CNR2X1 U1052 ( .A(n38), .B(n52), .Z(n837) );
  CNR2X1 U1053 ( .A(n912), .B(n911), .Z(n795) );
  CNR2X1 U1054 ( .A(n52), .B(n16), .Z(n755) );
  CNR2X1 U1055 ( .A(n42), .B(n21), .Z(n695) );
  CNR2X1 U1056 ( .A(n48), .B(n910), .Z(n786) );
  CNR2X1 U1057 ( .A(n912), .B(n52), .Z(n809) );
  CNR2X1 U1058 ( .A(n40), .B(n18), .Z(n732) );
  CNR2X1 U1059 ( .A(n40), .B(n44), .Z(n866) );
  CNR2X1 U1060 ( .A(n38), .B(n46), .Z(n861) );
  CNR2X1 U1061 ( .A(n38), .B(n48), .Z(n854) );
  CNR2X1 U1062 ( .A(n911), .B(n15), .Z(n767) );
  CNR2X1 U1063 ( .A(n48), .B(n20), .Z(n703) );
  CNR2X1 U1064 ( .A(n34), .B(n27), .Z(n654) );
  CNR2X1 U1065 ( .A(n38), .B(n19), .Z(n720) );
  CNR2X1 U1066 ( .A(n34), .B(n21), .Z(n699) );
  CNR2X1 U1067 ( .A(n38), .B(n42), .Z(n872) );
  CEOXL U1068 ( .A(n61), .B(n96), .Z(product[26]) );
  CND2X1 U1069 ( .A(n216), .B(n95), .Z(n61) );
  CNR2X1 U1070 ( .A(n912), .B(n16), .Z(n753) );
  CNR2X1 U1071 ( .A(n44), .B(n22), .Z(n684) );
  CNR2X1 U1072 ( .A(n32), .B(n23), .Z(n681) );
  CNR2X1 U1073 ( .A(n48), .B(n912), .Z(n811) );
  CNR2X1 U1074 ( .A(n36), .B(n18), .Z(n734) );
  CNR2X1 U1075 ( .A(n34), .B(n19), .Z(n722) );
  CNR2X1 U1076 ( .A(n32), .B(n24), .Z(n673) );
  CNR2X1 U1077 ( .A(n44), .B(n50), .Z(n843) );
  CNR2X1 U1078 ( .A(n40), .B(n15), .Z(n776) );
  CNR2X1 U1079 ( .A(n36), .B(n17), .Z(n748) );
  CNR2X1 U1080 ( .A(n910), .B(n42), .Z(n789) );
  CNR2X1 U1081 ( .A(n32), .B(n28), .Z(n651) );
  COR2X1 U1082 ( .A(n645), .B(n882), .Z(n1003) );
  CNR2X1 U1083 ( .A(n50), .B(n911), .Z(n798) );
  CAOR1X1 U1084 ( .A(n1005), .B(n93), .C(n90), .Z(n1004) );
  CNR2X1 U1085 ( .A(n38), .B(n24), .Z(n670) );
  CNR2X1 U1086 ( .A(n44), .B(n912), .Z(n813) );
  CNR2X1 U1087 ( .A(n38), .B(n15), .Z(n777) );
  CNR2X1 U1088 ( .A(n40), .B(n50), .Z(n845) );
  CNR2X1 U1089 ( .A(n38), .B(n23), .Z(n678) );
  CNR2X1 U1090 ( .A(n32), .B(n19), .Z(n723) );
  CNR2X1 U1091 ( .A(n38), .B(n16), .Z(n762) );
  CNR2X1 U1092 ( .A(n38), .B(n50), .Z(n846) );
  CNR2X1 U1093 ( .A(n32), .B(n46), .Z(n864) );
  CNR2X1 U1094 ( .A(n48), .B(n15), .Z(n772) );
  CNR2X1 U1095 ( .A(n54), .B(n15), .Z(n769) );
  CNR2X1 U1096 ( .A(n32), .B(n26), .Z(n660) );
  CNR2X1 U1097 ( .A(n44), .B(n20), .Z(n705) );
  CNR2X1 U1098 ( .A(n46), .B(n911), .Z(n800) );
  CNR2X1 U1099 ( .A(n44), .B(n910), .Z(n788) );
  CNR2X1 U1100 ( .A(n40), .B(n16), .Z(n761) );
  CNR2X1 U1101 ( .A(n50), .B(n20), .Z(n702) );
  CNR2X1 U1102 ( .A(n32), .B(n29), .Z(n648) );
  CNR2X1 U1103 ( .A(n50), .B(n15), .Z(n771) );
  CNR2X1 U1104 ( .A(n44), .B(n16), .Z(n759) );
  CNR2X1 U1105 ( .A(n46), .B(n15), .Z(n773) );
  CNR2X1 U1106 ( .A(n42), .B(n17), .Z(n745) );
  CNR2X1 U1107 ( .A(n54), .B(n911), .Z(n796) );
  CNR2X1 U1108 ( .A(n40), .B(n20), .Z(n707) );
  CEOX1 U1109 ( .A(n646), .B(n647), .Z(n253) );
  CND2X1 U1110 ( .A(n645), .B(n882), .Z(n209) );
  CND2X1 U1111 ( .A(n639), .B(n641), .Z(n201) );
  CND2X1 U1112 ( .A(n335), .B(n358), .Z(n92) );
  CNR2X1 U1113 ( .A(n44), .B(n23), .Z(n675) );
  CND2X1 U1114 ( .A(n643), .B(n644), .Z(n204) );
  COR2X1 U1115 ( .A(n335), .B(n358), .Z(n1005) );
  COR2X1 U1116 ( .A(n639), .B(n641), .Z(n1006) );
  CEOXL U1117 ( .A(n63), .B(n104), .Z(product[24]) );
  CND2X1 U1118 ( .A(n218), .B(n103), .Z(n63) );
  CNR2XL U1119 ( .A(n1050), .B(n1048), .Z(n105) );
  COND1XL U1120 ( .A(n1047), .B(n1050), .C(n1049), .Z(n106) );
  CIVX4 U1121 ( .A(b[1]), .Z(n34) );
  CND2XL U1122 ( .A(n1055), .B(n1054), .Z(n147) );
  CANR1XL U1123 ( .A(n155), .B(n1055), .C(n150), .Z(n148) );
  CND2XL U1124 ( .A(n221), .B(n1057), .Z(n114) );
  CANR1XL U1125 ( .A(n122), .B(n221), .C(n117), .Z(n115) );
  CANR1XL U1126 ( .A(n142), .B(n1056), .C(n135), .Z(n133) );
  CIVX2 U1127 ( .A(b[21]), .Z(n21) );
  CIVX2 U1128 ( .A(b[14]), .Z(n910) );
  CIVX2 U1129 ( .A(b[16]), .Z(n16) );
  CNR2X1 U1130 ( .A(n1009), .B(n1008), .Z(n102) );
  CNR2X1 U1131 ( .A(n359), .B(n1013), .Z(n94) );
  CIVX2 U1132 ( .A(b[18]), .Z(n18) );
  CNR2XL U1133 ( .A(n38), .B(n20), .Z(n708) );
  CNR2XL U1134 ( .A(n32), .B(n42), .Z(n875) );
  CNR2XL U1135 ( .A(n34), .B(n52), .Z(n839) );
  CIVX2 U1136 ( .A(b[19]), .Z(n19) );
  CIVX2 U1137 ( .A(b[20]), .Z(n20) );
  COR2X1 U1138 ( .A(n1012), .B(n1010), .Z(n1007) );
  CNR2X1 U1139 ( .A(n34), .B(n20), .Z(n710) );
  CNR2XL U1140 ( .A(n40), .B(n25), .Z(n662) );
  CNR2X1 U1141 ( .A(n46), .B(n20), .Z(n704) );
  CNR2XL U1142 ( .A(n34), .B(n18), .Z(n735) );
  CNR2XL U1143 ( .A(n48), .B(n42), .Z(n852) );
  CNR2XL U1144 ( .A(n32), .B(n25), .Z(n666) );
  CNR2XL U1145 ( .A(n36), .B(n42), .Z(n873) );
  CNR2XL U1146 ( .A(n32), .B(n15), .Z(n780) );
  CND2X1 U1147 ( .A(n1012), .B(n1010), .Z(n100) );
  CND2X1 U1148 ( .A(n1009), .B(n1008), .Z(n103) );
  CND2X1 U1149 ( .A(n359), .B(n1013), .Z(n95) );
  CEOX1 U1150 ( .A(n71), .B(n153), .Z(product[16]) );
  CND2XL U1151 ( .A(n1055), .B(n1038), .Z(n71) );
  CANR1XL U1152 ( .A(n1054), .B(n158), .C(n155), .Z(n153) );
  CENX1 U1153 ( .A(n138), .B(n69), .Z(product[18]) );
  CND2XL U1154 ( .A(n1056), .B(n1041), .Z(n69) );
  COND1XL U1155 ( .A(n1040), .B(n145), .C(n1039), .Z(n138) );
  CENX1 U1156 ( .A(n131), .B(n68), .Z(product[19]) );
  CND2XL U1157 ( .A(n223), .B(n1042), .Z(n68) );
  COND1XL U1158 ( .A(n132), .B(n145), .C(n133), .Z(n131) );
  CENX1 U1159 ( .A(n109), .B(n64), .Z(product[23]) );
  CND2XL U1160 ( .A(n219), .B(n1049), .Z(n64) );
  COND1XL U1161 ( .A(n1048), .B(n112), .C(n1047), .Z(n109) );
  CENX1 U1162 ( .A(n1031), .B(n1051), .Z(n1091) );
  CENX1 U1163 ( .A(n164), .B(n1035), .Z(n1089) );
  COND1XL U1164 ( .A(n1034), .B(n167), .C(n1033), .Z(n164) );
  CENX1 U1165 ( .A(n158), .B(n72), .Z(product[15]) );
  CND2XL U1166 ( .A(n1054), .B(n1037), .Z(n72) );
  CENX1 U1167 ( .A(n125), .B(n67), .Z(product[20]) );
  CND2XL U1168 ( .A(n1057), .B(n1044), .Z(n67) );
  CEOX1 U1169 ( .A(n175), .B(n1032), .Z(n1090) );
  CANR1XL U1170 ( .A(n1053), .B(n1051), .C(n1052), .Z(n175) );
  CEOX1 U1171 ( .A(n74), .B(n167), .Z(product[13]) );
  CND2X1 U1172 ( .A(n229), .B(n1033), .Z(n74) );
  CEOX1 U1173 ( .A(n70), .B(n145), .Z(product[17]) );
  CND2XL U1174 ( .A(n225), .B(n1039), .Z(n70) );
  CEOX1 U1175 ( .A(n66), .B(n120), .Z(product[21]) );
  CND2XL U1176 ( .A(n221), .B(n1045), .Z(n66) );
  CANR1XL U1177 ( .A(n1057), .B(n125), .C(n122), .Z(n120) );
  CEOX1 U1178 ( .A(n65), .B(n112), .Z(product[22]) );
  CNR2XL U1179 ( .A(n885), .B(a[1]), .Z(n212) );
  CIVX2 U1180 ( .A(n84), .Z(product[2]) );
  CIVX2 U1181 ( .A(n100), .Z(n98) );
  CIVX2 U1182 ( .A(n92), .Z(n90) );
  CIVX2 U1183 ( .A(b[30]), .Z(n30) );
  CIVX2 U1184 ( .A(b[29]), .Z(n29) );
  CIVX2 U1185 ( .A(b[27]), .Z(n27) );
  CIVX2 U1186 ( .A(b[26]), .Z(n26) );
  CIVX2 U1187 ( .A(b[25]), .Z(n25) );
  CIVX2 U1188 ( .A(b[24]), .Z(n24) );
  CIVX2 U1189 ( .A(n203), .Z(n237) );
  CIVX2 U1190 ( .A(n195), .Z(n235) );
  CIVX2 U1191 ( .A(n187), .Z(n233) );
  CIVX2 U1192 ( .A(b[23]), .Z(n23) );
  CIVX2 U1193 ( .A(n1034), .Z(n229) );
  CIVX2 U1194 ( .A(n1043), .Z(n223) );
  CIVX2 U1195 ( .A(n1048), .Z(n220) );
  CIVX2 U1196 ( .A(n1050), .Z(n219) );
  CIVX2 U1197 ( .A(n102), .Z(n218) );
  CIVX2 U1198 ( .A(n94), .Z(n216) );
  CIVX2 U1199 ( .A(n209), .Z(n207) );
  CIVX2 U1200 ( .A(n201), .Z(n199) );
  CIVX2 U1201 ( .A(n193), .Z(n191) );
  CIVX2 U1202 ( .A(n185), .Z(n183) );
  CIVX2 U1203 ( .A(n174), .Z(n172) );
  CIVX2 U1204 ( .A(n1029), .Z(n167) );
  CIVX2 U1205 ( .A(n159), .Z(n158) );
  CIVX2 U1206 ( .A(n1037), .Z(n155) );
  CIVX2 U1207 ( .A(n146), .Z(n145) );
  CIVX2 U1208 ( .A(n1039), .Z(n142) );
  CIVX2 U1209 ( .A(n1040), .Z(n225) );
  CIVX2 U1210 ( .A(n1044), .Z(n122) );
  CIVX2 U1211 ( .A(n1045), .Z(n117) );
  CIVX2 U1212 ( .A(n1046), .Z(n221) );
  CIVX2 U1213 ( .A(n113), .Z(n112) );
endmodule


module calc_DW02_mult_2_stage_9 ( A, B, TC, CLK, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC, CLK;
  wire   n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, \B_extended[32] ,
         n6, n8, n10, n12, n14, n16, n18, n20, n22, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34;
  assign \B_extended[32]  = B[31];

  calc_DW_mult_tc_20 mult_96 ( .a({\B_extended[32] , A}), .b({\B_extended[32] , 
        \B_extended[32] , B[30:0]}), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, PRODUCT[31:11], n35, n36, n37, n38, n39, n40, 
        n41, n42, n43, SYNOPSYS_UNCONNECTED__34, n44}), .dw2_CLK(CLK) );
  CFD1QXL clk_r_REG56_S1 ( .D(n43), .CP(CLK), .Q(n26) );
  CFD1QXL clk_r_REG57_S1 ( .D(n42), .CP(CLK), .Q(n27) );
  CFD1QXL clk_r_REG52_S1 ( .D(n39), .CP(CLK), .Q(n30) );
  CFD1QXL clk_r_REG55_S1 ( .D(n40), .CP(CLK), .Q(n29) );
  CFD1QXL clk_r_REG54_S1 ( .D(n41), .CP(CLK), .Q(n28) );
  CFD1QXL clk_r_REG51_S1 ( .D(n36), .CP(CLK), .Q(n33) );
  CFD1QXL clk_r_REG50_S1 ( .D(n37), .CP(CLK), .Q(n32) );
  CFD1QXL clk_r_REG53_S1 ( .D(n38), .CP(CLK), .Q(n31) );
  CFD1QXL clk_r_REG45_S1 ( .D(n35), .CP(CLK), .Q(n34) );
  CFD1QXL clk_r_REG59_S1 ( .D(n44), .CP(CLK), .Q(n25) );
  CIVDXL U1 ( .A(n33), .Z1(n6) );
  CNIVX1 U2 ( .A(n6), .Z(PRODUCT[9]) );
  CIVDXL U3 ( .A(n29), .Z1(n8) );
  CNIVX1 U4 ( .A(n8), .Z(PRODUCT[5]) );
  CIVDXL U5 ( .A(n25), .Z1(n10) );
  CNIVX1 U6 ( .A(n10), .Z(PRODUCT[0]) );
  CIVDXL U7 ( .A(n26), .Z1(n12) );
  CNIVX1 U8 ( .A(n12), .Z(PRODUCT[2]) );
  CIVDXL U9 ( .A(n31), .Z1(n14) );
  CNIVX1 U10 ( .A(n14), .Z(PRODUCT[7]) );
  CIVDXL U11 ( .A(n27), .Z1(n16) );
  CNIVX1 U12 ( .A(n16), .Z(PRODUCT[3]) );
  CIVDXL U13 ( .A(n32), .Z1(n18) );
  CNIVX1 U14 ( .A(n18), .Z(PRODUCT[8]) );
  CIVDXL U15 ( .A(n28), .Z1(n20) );
  CNIVX1 U16 ( .A(n20), .Z(PRODUCT[4]) );
  CIVDXL U17 ( .A(n34), .Z1(n22) );
  CNIVX1 U18 ( .A(n22), .Z(PRODUCT[10]) );
  CIVDXL U19 ( .A(n30), .Z1(n24) );
  CNIVX1 U20 ( .A(n24), .Z(PRODUCT[6]) );
endmodule


module calc_DW_mult_tc_21 ( a, b, product, dw1_CLK );
  input [32:0] a;
  input [32:0] b;
  output [65:0] product;
  input dw1_CLK;
  wire   n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n32, n34, n36, n38, n40, n42, n44, n46, n48, n50, n52, n54,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n90, n92, n93, n94, n95, n96, n98, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n117,
         n118, n119, n120, n122, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n135, n137, n138, n139, n140, n142, n145, n146,
         n147, n148, n150, n152, n153, n155, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n172, n174,
         n175, n177, n179, n180, n181, n183, n185, n186, n187, n188, n189,
         n191, n193, n194, n195, n196, n197, n199, n201, n202, n203, n204,
         n205, n207, n209, n210, n212, n213, n216, n218, n219, n220, n221,
         n223, n225, n229, n233, n235, n237, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n885, n910, n911, n912, \b[0] , n1089, n1088, n1087, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056;
  assign product[0] = \b[0] ;
  assign \b[0]  = b[0];
  assign n1056 = dw1_CLK;

  CFA1X1 U50 ( .A(n282), .B(n86), .CI(n255), .CO(n85), .S(product[30]) );
  CFA1X1 U51 ( .A(n308), .B(n87), .CI(n283), .CO(n86), .S(product[29]) );
  CFA1X1 U52 ( .A(n334), .B(n1002), .CI(n309), .CO(n87), .S(product[28]) );
  CEO3X2 U257 ( .A(n260), .B(n243), .C(n242), .Z(n241) );
  CEO3X2 U258 ( .A(n245), .B(n262), .C(n244), .Z(n242) );
  CEO3X2 U259 ( .A(n246), .B(n247), .C(n264), .Z(n243) );
  CEO3X2 U260 ( .A(n248), .B(n268), .C(n266), .Z(n244) );
  CEO3X2 U261 ( .A(n249), .B(n250), .C(n270), .Z(n245) );
  CEO3X2 U262 ( .A(n274), .B(n251), .C(n252), .Z(n246) );
  CEO3X2 U263 ( .A(n276), .B(n272), .C(n253), .Z(n247) );
  CEO3X2 U266 ( .A(n667), .B(n674), .C(n682), .Z(n250) );
  CEO3X2 U268 ( .A(n701), .B(n649), .C(n751), .Z(n252) );
  CFA1X1 U270 ( .A(n1024), .B(n1025), .CI(n1023), .CO(n254), .S(n255) );
  CFA1X1 U271 ( .A(n288), .B(n286), .CI(n261), .CO(n256), .S(n257) );
  CFA1X1 U272 ( .A(n265), .B(n263), .CI(n290), .CO(n258), .S(n259) );
  CFA1X1 U273 ( .A(n269), .B(n267), .CI(n292), .CO(n260), .S(n261) );
  CFA1X1 U274 ( .A(n271), .B(n294), .CI(n296), .CO(n262), .S(n263) );
  CFA1X1 U275 ( .A(n275), .B(n277), .CI(n273), .CO(n264), .S(n265) );
  CFA1X1 U276 ( .A(n298), .B(n279), .CI(n300), .CO(n266), .S(n267) );
  CFA1X1 U277 ( .A(n281), .B(n302), .CI(n304), .CO(n268), .S(n269) );
  CFA1X1 U278 ( .A(n692), .B(n306), .CI(n713), .CO(n270), .S(n271) );
  CFA1X1 U279 ( .A(n725), .B(n683), .CI(n657), .CO(n272), .S(n273) );
  CFA1X1 U281 ( .A(n675), .B(n752), .CI(n650), .CO(n276), .S(n277) );
  CFA1X1 U282 ( .A(n702), .B(n766), .CI(n648), .CO(n278), .S(n279) );
  CHA1X1 U283 ( .A(a[15]), .B(n662), .CO(n280), .S(n281) );
  CFA1X1 U284 ( .A(n1021), .B(n1022), .CI(n1020), .CO(n282), .S(n283) );
  CFA1X1 U285 ( .A(n291), .B(n312), .CI(n289), .CO(n284), .S(n285) );
  CFA1X1 U286 ( .A(n316), .B(n314), .CI(n293), .CO(n286), .S(n287) );
  CFA1X1 U287 ( .A(n297), .B(n295), .CI(n318), .CO(n288), .S(n289) );
  CFA1X1 U288 ( .A(n301), .B(n320), .CI(n299), .CO(n290), .S(n291) );
  CFA1X1 U289 ( .A(n305), .B(n322), .CI(n303), .CO(n292), .S(n293) );
  CFA1X1 U290 ( .A(n328), .B(n326), .CI(n324), .CO(n294), .S(n295) );
  CFA1X1 U291 ( .A(n332), .B(n330), .CI(n307), .CO(n296), .S(n297) );
  CFA1X1 U292 ( .A(n714), .B(n693), .CI(n676), .CO(n298), .S(n299) );
  CFA1X1 U294 ( .A(n684), .B(n739), .CI(n753), .CO(n302), .S(n303) );
  CFA1X1 U295 ( .A(n703), .B(n654), .CI(n767), .CO(n304), .S(n305) );
  CHA1X1 U296 ( .A(n663), .B(n651), .CO(n306), .S(n307) );
  CFA1X1 U297 ( .A(n1018), .B(n1019), .CI(n1017), .CO(n308), .S(n309) );
  CFA1X1 U298 ( .A(n340), .B(n338), .CI(n315), .CO(n310), .S(n311) );
  CFA1X1 U299 ( .A(n342), .B(n317), .CI(n319), .CO(n312), .S(n313) );
  CFA1X1 U300 ( .A(n346), .B(n321), .CI(n344), .CO(n314), .S(n315) );
  CFA1X1 U301 ( .A(n331), .B(n323), .CI(n329), .CO(n316), .S(n317) );
  CFA1X1 U302 ( .A(n348), .B(n325), .CI(n327), .CO(n318), .S(n319) );
  CFA1X1 U303 ( .A(n354), .B(n352), .CI(n350), .CO(n320), .S(n321) );
  CFA1X1 U304 ( .A(n715), .B(n333), .CI(n356), .CO(n322), .S(n323) );
  CFA1X1 U305 ( .A(n727), .B(n694), .CI(n677), .CO(n324), .S(n325) );
  CFA1X1 U306 ( .A(n670), .B(n659), .CI(n740), .CO(n326), .S(n327) );
  CFA1X1 U307 ( .A(n685), .B(n754), .CI(n655), .CO(n328), .S(n329) );
  CFA1X1 U308 ( .A(n664), .B(n781), .CI(n768), .CO(n330), .S(n331) );
  CHA1X1 U309 ( .A(a[14]), .B(n704), .CO(n332), .S(n333) );
  CFA1X1 U310 ( .A(n1015), .B(n1016), .CI(n1014), .CO(n334), .S(n335) );
  CFA1X1 U311 ( .A(n364), .B(n362), .CI(n341), .CO(n336), .S(n337) );
  CFA1X1 U312 ( .A(n366), .B(n343), .CI(n345), .CO(n338), .S(n339) );
  CFA1X1 U313 ( .A(n370), .B(n347), .CI(n368), .CO(n340), .S(n341) );
  CFA1X1 U314 ( .A(n353), .B(n349), .CI(n351), .CO(n342), .S(n343) );
  CFA1X1 U315 ( .A(n374), .B(n355), .CI(n372), .CO(n344), .S(n345) );
  CFA1X1 U316 ( .A(n357), .B(n376), .CI(n378), .CO(n346), .S(n347) );
  CFA1X1 U317 ( .A(n741), .B(n380), .CI(n728), .CO(n348), .S(n349) );
  CFA1X1 U318 ( .A(n755), .B(n716), .CI(n695), .CO(n350), .S(n351) );
  CFA1X1 U320 ( .A(n705), .B(n660), .CI(n769), .CO(n354), .S(n355) );
  CHA1X1 U321 ( .A(n665), .B(n782), .CO(n356), .S(n357) );
  CFA1X1 U322 ( .A(n1012), .B(n1013), .CI(n1009), .CO(n358), .S(n359) );
  CFA1X1 U323 ( .A(n388), .B(n386), .CI(n365), .CO(n360), .S(n361) );
  CFA1X1 U324 ( .A(n390), .B(n367), .CI(n369), .CO(n362), .S(n363) );
  CFA1X1 U325 ( .A(n394), .B(n371), .CI(n392), .CO(n364), .S(n365) );
  CFA1X1 U326 ( .A(n373), .B(n375), .CI(n377), .CO(n366), .S(n367) );
  CFA1X1 U327 ( .A(n398), .B(n379), .CI(n396), .CO(n368), .S(n369) );
  CFA1X1 U328 ( .A(n402), .B(n400), .CI(n381), .CO(n370), .S(n371) );
  CFA1X1 U329 ( .A(n756), .B(n742), .CI(n729), .CO(n372), .S(n373) );
  CFA1X1 U330 ( .A(n770), .B(n717), .CI(n687), .CO(n374), .S(n375) );
  CFA1X1 U331 ( .A(n696), .B(n679), .CI(n672), .CO(n376), .S(n377) );
  CFA1X1 U332 ( .A(n706), .B(n783), .CI(n795), .CO(n378), .S(n379) );
  CHA1X1 U333 ( .A(a[13]), .B(n666), .CO(n380), .S(n381) );
  CFA1X1 U334 ( .A(n387), .B(n385), .CI(n406), .CO(n382), .S(n383) );
  CFA1X1 U335 ( .A(n391), .B(n389), .CI(n408), .CO(n384), .S(n385) );
  CFA1X1 U336 ( .A(n412), .B(n410), .CI(n393), .CO(n386), .S(n387) );
  CFA1X1 U337 ( .A(n397), .B(n395), .CI(n414), .CO(n388), .S(n389) );
  CFA1X1 U338 ( .A(n416), .B(n399), .CI(n401), .CO(n390), .S(n391) );
  CFA1X1 U339 ( .A(n422), .B(n420), .CI(n418), .CO(n392), .S(n393) );
  CFA1X1 U340 ( .A(n743), .B(n403), .CI(n424), .CO(n394), .S(n395) );
  CFA1X1 U341 ( .A(n757), .B(n697), .CI(n688), .CO(n396), .S(n397) );
  CFA1X1 U342 ( .A(n730), .B(n771), .CI(n784), .CO(n398), .S(n399) );
  CFA1X1 U343 ( .A(n718), .B(n680), .CI(n673), .CO(n400), .S(n401) );
  CHA1X1 U344 ( .A(n707), .B(n796), .CO(n402), .S(n403) );
  CFA1X1 U345 ( .A(n409), .B(n407), .CI(n428), .CO(n404), .S(n405) );
  CFA1X1 U346 ( .A(n413), .B(n430), .CI(n411), .CO(n406), .S(n407) );
  CFA1X1 U347 ( .A(n434), .B(n432), .CI(n415), .CO(n408), .S(n409) );
  CFA1X1 U348 ( .A(n423), .B(n436), .CI(n417), .CO(n410), .S(n411) );
  CFA1X1 U349 ( .A(n438), .B(n421), .CI(n419), .CO(n412), .S(n413) );
  CFA1X1 U350 ( .A(n425), .B(n440), .CI(n442), .CO(n414), .S(n415) );
  CFA1X1 U351 ( .A(n731), .B(n444), .CI(n719), .CO(n416), .S(n417) );
  CFA1X1 U352 ( .A(n758), .B(n689), .CI(n681), .CO(n418), .S(n419) );
  CFA1X1 U353 ( .A(n698), .B(n772), .CI(n797), .CO(n420), .S(n421) );
  CFA1X1 U354 ( .A(n744), .B(n785), .CI(n808), .CO(n422), .S(n423) );
  CHA1X1 U355 ( .A(a[12]), .B(n708), .CO(n424), .S(n425) );
  CFA1X1 U356 ( .A(n431), .B(n429), .CI(n448), .CO(n426), .S(n427) );
  CFA1X1 U357 ( .A(n435), .B(n450), .CI(n433), .CO(n428), .S(n429) );
  CFA1X1 U358 ( .A(n454), .B(n452), .CI(n437), .CO(n430), .S(n431) );
  CFA1X1 U359 ( .A(n443), .B(n456), .CI(n441), .CO(n432), .S(n433) );
  CFA1X1 U360 ( .A(n460), .B(n439), .CI(n458), .CO(n434), .S(n435) );
  CFA1X1 U361 ( .A(n464), .B(n462), .CI(n445), .CO(n436), .S(n437) );
  CFA1X1 U362 ( .A(n773), .B(n759), .CI(n745), .CO(n438), .S(n439) );
  CFA1X1 U363 ( .A(n720), .B(n699), .CI(n690), .CO(n440), .S(n441) );
  CFA1X1 U364 ( .A(n732), .B(n786), .CI(n809), .CO(n442), .S(n443) );
  CHA1X1 U365 ( .A(n709), .B(n798), .CO(n444), .S(n445) );
  CFA1X1 U366 ( .A(n451), .B(n449), .CI(n468), .CO(n446), .S(n447) );
  CFA1X1 U367 ( .A(n455), .B(n470), .CI(n453), .CO(n448), .S(n449) );
  CFA1X1 U368 ( .A(n457), .B(n472), .CI(n474), .CO(n450), .S(n451) );
  CFA1X1 U369 ( .A(n459), .B(n461), .CI(n463), .CO(n452), .S(n453) );
  CFA1X1 U370 ( .A(n480), .B(n476), .CI(n478), .CO(n454), .S(n455) );
  CFA1X1 U371 ( .A(n746), .B(n465), .CI(n482), .CO(n456), .S(n457) );
  CFA1X1 U372 ( .A(n760), .B(n721), .CI(n700), .CO(n458), .S(n459) );
  CFA1X1 U373 ( .A(n733), .B(n787), .CI(n774), .CO(n460), .S(n461) );
  CFA1X1 U374 ( .A(n820), .B(n799), .CI(n810), .CO(n462), .S(n463) );
  CHA1X1 U375 ( .A(a[11]), .B(n710), .CO(n464), .S(n465) );
  CFA1X1 U376 ( .A(n471), .B(n469), .CI(n486), .CO(n466), .S(n467) );
  CFA1X1 U377 ( .A(n490), .B(n488), .CI(n473), .CO(n468), .S(n469) );
  CFA1X1 U378 ( .A(n477), .B(n475), .CI(n492), .CO(n470), .S(n471) );
  CFA1X1 U379 ( .A(n494), .B(n481), .CI(n479), .CO(n472), .S(n473) );
  CFA1X1 U380 ( .A(n483), .B(n496), .CI(n498), .CO(n474), .S(n475) );
  CFA1X1 U381 ( .A(n775), .B(n500), .CI(n747), .CO(n476), .S(n477) );
  CFA1X1 U382 ( .A(n734), .B(n811), .CI(n722), .CO(n478), .S(n479) );
  CFA1X1 U383 ( .A(n761), .B(n800), .CI(n788), .CO(n480), .S(n481) );
  CHA1X1 U384 ( .A(n711), .B(n821), .CO(n482), .S(n483) );
  CFA1X1 U385 ( .A(n489), .B(n487), .CI(n504), .CO(n484), .S(n485) );
  CFA1X1 U386 ( .A(n493), .B(n506), .CI(n491), .CO(n486), .S(n487) );
  CFA1X1 U387 ( .A(n499), .B(n508), .CI(n510), .CO(n488), .S(n489) );
  CFA1X1 U388 ( .A(n512), .B(n497), .CI(n495), .CO(n490), .S(n491) );
  CFA1X1 U389 ( .A(n516), .B(n514), .CI(n501), .CO(n492), .S(n493) );
  CFA1X1 U390 ( .A(n789), .B(n776), .CI(n748), .CO(n494), .S(n495) );
  CFA1X1 U391 ( .A(n762), .B(n822), .CI(n723), .CO(n496), .S(n497) );
  CFA1X1 U392 ( .A(n831), .B(n801), .CI(n812), .CO(n498), .S(n499) );
  CHA1X1 U393 ( .A(a[10]), .B(n735), .CO(n500), .S(n501) );
  CFA1X1 U394 ( .A(n507), .B(n505), .CI(n520), .CO(n502), .S(n503) );
  CFA1X1 U395 ( .A(n511), .B(n509), .CI(n522), .CO(n504), .S(n505) );
  CFA1X1 U396 ( .A(n513), .B(n524), .CI(n515), .CO(n506), .S(n507) );
  CFA1X1 U397 ( .A(n530), .B(n526), .CI(n528), .CO(n508), .S(n509) );
  CFA1X1 U398 ( .A(n832), .B(n517), .CI(n532), .CO(n510), .S(n511) );
  CFA1X1 U400 ( .A(n777), .B(n823), .CI(n813), .CO(n514), .S(n515) );
  CHA1X1 U401 ( .A(n736), .B(n790), .CO(n516), .S(n517) );
  CFA1X1 U402 ( .A(n523), .B(n521), .CI(n536), .CO(n518), .S(n519) );
  CFA1X1 U403 ( .A(n540), .B(n538), .CI(n525), .CO(n520), .S(n521) );
  CFA1X1 U404 ( .A(n529), .B(n527), .CI(n531), .CO(n522), .S(n523) );
  CFA1X1 U405 ( .A(n533), .B(n542), .CI(n544), .CO(n524), .S(n525) );
  CFA1X1 U406 ( .A(n833), .B(n546), .CI(n764), .CO(n526), .S(n527) );
  CFA1X1 U407 ( .A(n778), .B(n791), .CI(n824), .CO(n528), .S(n529) );
  CFA1X1 U408 ( .A(n814), .B(n841), .CI(n803), .CO(n530), .S(n531) );
  CHA1X1 U409 ( .A(a[9]), .B(n750), .CO(n532), .S(n533) );
  CFA1X1 U410 ( .A(n539), .B(n537), .CI(n550), .CO(n534), .S(n535) );
  CFA1X1 U411 ( .A(n554), .B(n552), .CI(n541), .CO(n536), .S(n537) );
  CFA1X1 U412 ( .A(n556), .B(n545), .CI(n543), .CO(n538), .S(n539) );
  CFA1X1 U413 ( .A(n560), .B(n558), .CI(n547), .CO(n540), .S(n541) );
  CFA1X1 U414 ( .A(n825), .B(n804), .CI(n765), .CO(n542), .S(n543) );
  CFA1X1 U415 ( .A(n834), .B(n792), .CI(n842), .CO(n544), .S(n545) );
  CHA1X1 U416 ( .A(n779), .B(n815), .CO(n546), .S(n547) );
  CFA1X1 U417 ( .A(n553), .B(n551), .CI(n564), .CO(n548), .S(n549) );
  CFA1X1 U418 ( .A(n557), .B(n566), .CI(n555), .CO(n550), .S(n551) );
  CFA1X1 U419 ( .A(n570), .B(n559), .CI(n568), .CO(n552), .S(n553) );
  CFA1X1 U420 ( .A(n843), .B(n561), .CI(n572), .CO(n554), .S(n555) );
  CFA1X1 U421 ( .A(n816), .B(n826), .CI(n850), .CO(n556), .S(n557) );
  CFA1X1 U422 ( .A(n835), .B(n805), .CI(n793), .CO(n558), .S(n559) );
  CHA1X1 U423 ( .A(a[8]), .B(n780), .CO(n560), .S(n561) );
  CFA1X1 U424 ( .A(n567), .B(n565), .CI(n576), .CO(n562), .S(n563) );
  CFA1X1 U425 ( .A(n571), .B(n578), .CI(n569), .CO(n564), .S(n565) );
  CFA1X1 U426 ( .A(n573), .B(n580), .CI(n582), .CO(n566), .S(n567) );
  CFA1X1 U427 ( .A(n817), .B(n584), .CI(n806), .CO(n568), .S(n569) );
  CFA1X1 U428 ( .A(n836), .B(n827), .CI(n851), .CO(n570), .S(n571) );
  CHA1X1 U429 ( .A(n844), .B(n794), .CO(n572), .S(n573) );
  CFA1X1 U430 ( .A(n579), .B(n577), .CI(n588), .CO(n574), .S(n575) );
  CFA1X1 U431 ( .A(n583), .B(n590), .CI(n581), .CO(n576), .S(n577) );
  CFA1X1 U432 ( .A(n594), .B(n592), .CI(n585), .CO(n578), .S(n579) );
  CFA1X1 U433 ( .A(n845), .B(n828), .CI(n818), .CO(n580), .S(n581) );
  CFA1X1 U434 ( .A(n837), .B(n858), .CI(n807), .CO(n582), .S(n583) );
  CHA1X1 U435 ( .A(a[7]), .B(n852), .CO(n584), .S(n585) );
  CFA1X1 U436 ( .A(n591), .B(n589), .CI(n598), .CO(n586), .S(n587) );
  CFA1X1 U437 ( .A(n602), .B(n593), .CI(n600), .CO(n588), .S(n589) );
  CFA1X1 U438 ( .A(n846), .B(n595), .CI(n604), .CO(n590), .S(n591) );
  CFA1X1 U439 ( .A(n859), .B(n829), .CI(n853), .CO(n592), .S(n593) );
  CHA1X1 U440 ( .A(n838), .B(n819), .CO(n594), .S(n595) );
  CFA1X1 U441 ( .A(n601), .B(n599), .CI(n608), .CO(n596), .S(n597) );
  CFA1X1 U442 ( .A(n605), .B(n603), .CI(n610), .CO(n598), .S(n599) );
  CFA1X1 U443 ( .A(n854), .B(n612), .CI(n847), .CO(n600), .S(n601) );
  CFA1X1 U444 ( .A(n865), .B(n860), .CI(n830), .CO(n602), .S(n603) );
  CHA1X1 U445 ( .A(a[6]), .B(n839), .CO(n604), .S(n605) );
  CFA1X1 U446 ( .A(n611), .B(n609), .CI(n616), .CO(n606), .S(n607) );
  CFA1X1 U447 ( .A(n620), .B(n618), .CI(n613), .CO(n608), .S(n609) );
  CFA1X1 U448 ( .A(n855), .B(n866), .CI(n861), .CO(n610), .S(n611) );
  CHA1X1 U449 ( .A(n840), .B(n848), .CO(n612), .S(n613) );
  CFA1X1 U450 ( .A(n624), .B(n617), .CI(n619), .CO(n614), .S(n615) );
  CFA1X1 U451 ( .A(n862), .B(n621), .CI(n626), .CO(n616), .S(n617) );
  CFA1X1 U452 ( .A(n867), .B(n856), .CI(n849), .CO(n618), .S(n619) );
  CHA1X1 U453 ( .A(a[5]), .B(n871), .CO(n620), .S(n621) );
  CFA1X1 U454 ( .A(n627), .B(n625), .CI(n630), .CO(n622), .S(n623) );
  CFA1X1 U455 ( .A(n868), .B(n632), .CI(n863), .CO(n624), .S(n625) );
  CHA1X1 U456 ( .A(n872), .B(n857), .CO(n626), .S(n627) );
  CFA1X1 U457 ( .A(n636), .B(n631), .CI(n633), .CO(n628), .S(n629) );
  CFA1X1 U458 ( .A(n876), .B(n869), .CI(n864), .CO(n630), .S(n631) );
  CHA1X1 U459 ( .A(a[4]), .B(n873), .CO(n632), .S(n633) );
  CFA1X1 U460 ( .A(n877), .B(n637), .CI(n640), .CO(n634), .S(n635) );
  CHA1X1 U461 ( .A(n874), .B(n870), .CO(n636), .S(n637) );
  CHA1X1 U463 ( .A(a[3]), .B(n875), .CO(n640), .S(n641) );
  CHA1X1 U464 ( .A(n881), .B(n879), .CO(n642), .S(n643) );
  CFD1QXL clk_r_REG49_S1 ( .D(n995), .CP(n1056), .Q(n1051) );
  CFD1QXL clk_r_REG48_S1 ( .D(n177), .CP(n1056), .Q(n1050) );
  CFD1QXL clk_r_REG0_S1 ( .D(n257), .CP(n1056), .Q(n1025) );
  CFD1QXL clk_r_REG44_S1 ( .D(n165), .CP(n1056), .Q(n1032) );
  CFD1QXL clk_r_REG43_S1 ( .D(n166), .CP(n1056), .Q(n1031) );
  CFD1QXL clk_r_REG6_S1 ( .D(n259), .CP(n1056), .Q(n1024) );
  CFD1QXL clk_r_REG36_S1 ( .D(n73), .CP(n1056), .Q(n1033) );
  CFD1QXL clk_r_REG41_S1 ( .D(n75), .CP(n1056), .Q(n1030) );
  CFD1QXL clk_r_REG47_S1 ( .D(n76), .CP(n1056), .Q(n1029) );
  CFD1QXL clk_r_REG1_S1 ( .D(n240), .CP(n1056), .Q(n1026) );
  CFD1QXL clk_r_REG46_S1 ( .D(n180), .CP(n1056), .Q(n1049) );
  CFD1QXL clk_r_REG38_S1 ( .D(n160), .CP(n1056), .Q(n1034) );
  CFD1QXL clk_r_REG37_S1 ( .D(n161), .CP(n1056), .Q(n1028) );
  CFD1QXL clk_r_REG4_S1 ( .D(n285), .CP(n1056), .Q(n1022) );
  CFD1QXL clk_r_REG42_S1 ( .D(n168), .CP(n1056), .Q(n1027) );
  CFD1QXL clk_r_REG35_S1 ( .D(n139), .CP(n1056), .Q(n1038) );
  CFD1QXL clk_r_REG21_S1 ( .D(n108), .CP(n1056), .Q(n1047) );
  CFD1QXL clk_r_REG11_S1 ( .D(n310), .CP(n1056), .Q(n1020) );
  CFD1QXL clk_r_REG9_S1 ( .D(n336), .CP(n1056), .Q(n1017) );
  CFD1QXL clk_r_REG7_S1 ( .D(n360), .CP(n1056), .Q(n1014) );
  CFD1QXL clk_r_REG16_S1 ( .D(n384), .CP(n1056), .Q(n1009) );
  CFD1QXL clk_r_REG5_S1 ( .D(n287), .CP(n1056), .Q(n1021) );
  CFD1QXL clk_r_REG2_S1 ( .D(n313), .CP(n1056), .Q(n1018) );
  CFD1QXL clk_r_REG13_S1 ( .D(n339), .CP(n1056), .Q(n1015) );
  CFD1QXL clk_r_REG58_S1 ( .D(n363), .CP(n1056), .Q(n1012) );
  CFD1QXL clk_r_REG26_S1 ( .D(n119), .CP(n1056), .Q(n1043) );
  CFD1QXL clk_r_REG24_S1 ( .D(n124), .CP(n1056), .Q(n1042) );
  CFD1QXL clk_r_REG32_S1 ( .D(n152), .CP(n1056), .Q(n1036) );
  CFD1QXL clk_r_REG28_S1 ( .D(n137), .CP(n1056), .Q(n1039) );
  CFD1QXL clk_r_REG39_S1 ( .D(n157), .CP(n1056), .Q(n1035) );
  CFD1QXL clk_r_REG15_S1 ( .D(n405), .CP(n1056), .Q(n1007) );
  CFD1QXL clk_r_REG19_S1 ( .D(n111), .CP(n1056), .Q(n1045) );
  CFD1QXL clk_r_REG17_S1 ( .D(n382), .CP(n1056), .Q(n1011) );
  CFD1QXL clk_r_REG14_S1 ( .D(n404), .CP(n1056), .Q(n1008) );
  CFD1QXL clk_r_REG23_S1 ( .D(n426), .CP(n1056), .Q(n1006) );
  CFD1QXL clk_r_REG22_S1 ( .D(n107), .CP(n1056), .Q(n1048) );
  CFD1QXL clk_r_REG33_S1 ( .D(n992), .CP(n1056), .Q(n1053) );
  CFD1QXL clk_r_REG29_S1 ( .D(n993), .CP(n1056), .Q(n1054) );
  CFD1QXL clk_r_REG20_S1 ( .D(n110), .CP(n1056), .Q(n1046) );
  CFD1QXL clk_r_REG34_S1 ( .D(n140), .CP(n1056), .Q(n1037) );
  CFD1QXL clk_r_REG25_S1 ( .D(n994), .CP(n1056), .Q(n1055) );
  CFD1QXL clk_r_REG40_S1 ( .D(n998), .CP(n1056), .Q(n1052) );
  CFD1QXL clk_r_REG8_S1 ( .D(n361), .CP(n1056), .Q(n1013) );
  CFD1QXL clk_r_REG3_S1 ( .D(n284), .CP(n1056), .Q(n1023) );
  CFD1QXL clk_r_REG12_S1 ( .D(n311), .CP(n1056), .Q(n1019) );
  CFD1QXL clk_r_REG30_S1 ( .D(n130), .CP(n1056), .Q(n1040) );
  CFD1QXL clk_r_REG31_S1 ( .D(n129), .CP(n1056), .Q(n1041) );
  CFD1QXL clk_r_REG10_S1 ( .D(n337), .CP(n1056), .Q(n1016) );
  CFD1QXL clk_r_REG27_S1 ( .D(n118), .CP(n1056), .Q(n1044) );
  CFD1QX2 clk_r_REG18_S1 ( .D(n383), .CP(n1056), .Q(n1010) );
  CIVX1 U754 ( .A(b[24]), .Z(n24) );
  CNR2XL U755 ( .A(n32), .B(n48), .Z(n857) );
  CNR2XL U756 ( .A(n32), .B(n50), .Z(n849) );
  CNR2XL U757 ( .A(n32), .B(n38), .Z(n882) );
  CNR2XL U758 ( .A(n32), .B(n912), .Z(n819) );
  CNR2XL U759 ( .A(n32), .B(n911), .Z(n807) );
  CNR2XL U760 ( .A(n32), .B(n910), .Z(n794) );
  CNR2XL U761 ( .A(n32), .B(n27), .Z(n655) );
  CIVX4 U762 ( .A(b[17]), .Z(n17) );
  COND1X1 U763 ( .A(n1041), .B(n133), .C(n1040), .Z(n128) );
  CIVXL U764 ( .A(n126), .Z(n125) );
  CNR2X1 U765 ( .A(n32), .B(n20), .Z(n711) );
  CNR2X1 U766 ( .A(n32), .B(n17), .Z(n750) );
  CNR2IX1 U767 ( .B(a[1]), .A(n17), .Z(n749) );
  CNR2X1 U768 ( .A(n54), .B(n17), .Z(n739) );
  CNR2X1 U769 ( .A(n44), .B(n17), .Z(n744) );
  CNR2X2 U770 ( .A(n42), .B(n17), .Z(n745) );
  CIVX8 U771 ( .A(\b[0] ), .Z(n32) );
  CFA1XL U772 ( .A(n668), .B(n653), .CI(n738), .CO(n274), .S(n275) );
  CEO3X1 U773 ( .A(n258), .B(n241), .C(n256), .Z(n240) );
  CNIVX1 U774 ( .A(n1089), .Z(product[11]) );
  CNIVX1 U775 ( .A(n1088), .Z(product[12]) );
  CNIVX1 U776 ( .A(n1087), .Z(product[14]) );
  CFA1XL U777 ( .A(n749), .B(n802), .CI(n990), .CO(n512), .S(n513) );
  COND1X2 U778 ( .A(n94), .B(n96), .C(n95), .Z(n93) );
  CANR1X2 U779 ( .A(n1005), .B(n101), .C(n98), .Z(n96) );
  CIVX1 U780 ( .A(n1036), .Z(n150) );
  COND1X2 U781 ( .A(n102), .B(n104), .C(n103), .Z(n101) );
  CANR1X2 U782 ( .A(n105), .B(n113), .C(n106), .Z(n104) );
  CHA1XL U783 ( .A(a[2]), .B(n883), .CO(n644), .S(n645) );
  CIVX4 U784 ( .A(b[2]), .Z(n36) );
  CFA1XL U785 ( .A(n726), .B(n669), .CI(n658), .CO(n300), .S(n301) );
  CNR2X1 U786 ( .A(n36), .B(n26), .Z(n658) );
  CFA1XL U787 ( .A(n686), .B(n678), .CI(n671), .CO(n352), .S(n353) );
  CIVXL U788 ( .A(n763), .Z(n989) );
  CIVX2 U789 ( .A(n989), .Z(n990) );
  CNR2XL U790 ( .A(n36), .B(n46), .Z(n862) );
  CNR2XL U791 ( .A(n36), .B(n50), .Z(n847) );
  CNR2XL U792 ( .A(n36), .B(n40), .Z(n877) );
  CNR2XL U793 ( .A(n36), .B(n52), .Z(n838) );
  CNR2XL U794 ( .A(n36), .B(n48), .Z(n855) );
  CNR2XL U795 ( .A(n36), .B(n28), .Z(n649) );
  CNR2XL U796 ( .A(n36), .B(n911), .Z(n805) );
  COR2XL U797 ( .A(n32), .B(n36), .Z(n1000) );
  CNR2XL U798 ( .A(n36), .B(n27), .Z(n653) );
  CNR2XL U799 ( .A(n36), .B(n24), .Z(n671) );
  CNR2XL U800 ( .A(n34), .B(n36), .Z(n883) );
  CNR2XL U801 ( .A(n36), .B(n16), .Z(n763) );
  CNR2XL U802 ( .A(n36), .B(n15), .Z(n778) );
  CNR2XL U803 ( .A(n36), .B(n910), .Z(n792) );
  CFA1XL U804 ( .A(n880), .B(n642), .CI(n878), .CO(n638), .S(n639) );
  CIVXL U805 ( .A(n181), .Z(n180) );
  CANR1X1 U806 ( .A(n997), .B(n186), .C(n183), .Z(n181) );
  COND1X1 U807 ( .A(n147), .B(n159), .C(n148), .Z(n146) );
  CANR1X1 U808 ( .A(n1034), .B(n1027), .C(n1028), .Z(n159) );
  COND1X2 U809 ( .A(n114), .B(n126), .C(n115), .Z(n113) );
  CANR1X2 U810 ( .A(n146), .B(n127), .C(n128), .Z(n126) );
  CNR2XL U811 ( .A(n36), .B(n25), .Z(n664) );
  CNR2XL U812 ( .A(n38), .B(n27), .Z(n652) );
  CNR2XL U813 ( .A(n50), .B(n19), .Z(n714) );
  CNR2XL U814 ( .A(n52), .B(n18), .Z(n726) );
  CNR2XL U815 ( .A(n42), .B(n25), .Z(n661) );
  CNR2XL U816 ( .A(n40), .B(n22), .Z(n686) );
  CNR2XL U817 ( .A(n912), .B(n17), .Z(n738) );
  CNR2X1 U818 ( .A(n38), .B(n40), .Z(n876) );
  CND2XL U819 ( .A(n1054), .B(n225), .Z(n132) );
  CEOXL U820 ( .A(n197), .B(n80), .Z(product[7]) );
  CANR1XL U821 ( .A(n210), .B(n1001), .C(n207), .Z(n205) );
  CNR2XL U822 ( .A(n42), .B(n52), .Z(n835) );
  CNR2XL U823 ( .A(n38), .B(n912), .Z(n816) );
  CNR2XL U824 ( .A(n912), .B(n15), .Z(n768) );
  CNR2XL U825 ( .A(n42), .B(n15), .Z(n775) );
  CNR2XL U826 ( .A(n40), .B(n52), .Z(n836) );
  CNR2XL U827 ( .A(n912), .B(n910), .Z(n782) );
  CNR2XL U828 ( .A(n36), .B(n912), .Z(n817) );
  CNR2X1 U829 ( .A(n34), .B(n23), .Z(n680) );
  CNR2XL U830 ( .A(n32), .B(n52), .Z(n840) );
  CNR2XL U831 ( .A(n38), .B(n44), .Z(n867) );
  CNR2XL U832 ( .A(n46), .B(n42), .Z(n859) );
  CNR2XL U833 ( .A(n32), .B(n40), .Z(n879) );
  CNR2XL U834 ( .A(n40), .B(n912), .Z(n815) );
  CNR2XL U835 ( .A(n32), .B(n28), .Z(n651) );
  CNR2XL U836 ( .A(n36), .B(n44), .Z(n868) );
  CNR2XL U837 ( .A(n46), .B(n52), .Z(n833) );
  CNR2XL U838 ( .A(n44), .B(n42), .Z(n865) );
  CNR2XL U839 ( .A(n32), .B(n44), .Z(n870) );
  CNR2XL U840 ( .A(n40), .B(n910), .Z(n790) );
  CNR2XL U841 ( .A(n32), .B(n30), .Z(n646) );
  CNR2XL U842 ( .A(n36), .B(n38), .Z(n880) );
  CIVX2 U843 ( .A(b[13]), .Z(n911) );
  CIVX2 U844 ( .A(b[14]), .Z(n910) );
  CIVX2 U845 ( .A(b[15]), .Z(n15) );
  CIVX3 U846 ( .A(b[10]), .Z(n52) );
  CIVX3 U847 ( .A(b[9]), .Z(n50) );
  CND2XL U848 ( .A(n885), .B(a[1]), .Z(n213) );
  CND2XL U849 ( .A(n997), .B(n185), .Z(n77) );
  CNR2XL U850 ( .A(n427), .B(n446), .Z(n107) );
  CNR2XL U851 ( .A(n447), .B(n466), .Z(n110) );
  CNR2XL U852 ( .A(n467), .B(n484), .Z(n118) );
  CNR2XL U853 ( .A(n162), .B(n165), .Z(n160) );
  CNR2XL U854 ( .A(n503), .B(n518), .Z(n129) );
  CNR2XL U855 ( .A(n535), .B(n548), .Z(n139) );
  CND2XL U856 ( .A(n485), .B(n502), .Z(n124) );
  CND2XL U857 ( .A(n503), .B(n518), .Z(n130) );
  CND2XL U858 ( .A(n996), .B(n174), .Z(n75) );
  CND2XL U859 ( .A(n535), .B(n548), .Z(n140) );
  CND2XL U860 ( .A(n995), .B(n179), .Z(n76) );
  CND2XL U861 ( .A(n549), .B(n562), .Z(n152) );
  CND2XL U862 ( .A(n519), .B(n534), .Z(n137) );
  CND2IXL U863 ( .B(n162), .A(n163), .Z(n73) );
  CIVXL U864 ( .A(n179), .Z(n177) );
  CND2XL U865 ( .A(n233), .B(n188), .Z(n78) );
  CND2XL U866 ( .A(n235), .B(n196), .Z(n80) );
  CND2XL U867 ( .A(n999), .B(n193), .Z(n79) );
  CND2XL U868 ( .A(n575), .B(n586), .Z(n163) );
  CND2XL U869 ( .A(n563), .B(n574), .Z(n157) );
  CANR1X1 U870 ( .A(n202), .B(n1004), .C(n199), .Z(n197) );
  CND2XL U871 ( .A(n237), .B(n204), .Z(n82) );
  CND2XL U872 ( .A(n1001), .B(n209), .Z(n83) );
  CND2XL U873 ( .A(n1004), .B(n201), .Z(n81) );
  CNR2XL U874 ( .A(n48), .B(n54), .Z(n822) );
  CNR2XL U875 ( .A(n34), .B(n44), .Z(n869) );
  CNR2XL U876 ( .A(n34), .B(n24), .Z(n672) );
  CNR2XL U877 ( .A(n36), .B(n23), .Z(n679) );
  CNR2XL U878 ( .A(n40), .B(n21), .Z(n696) );
  CNR2XL U879 ( .A(n46), .B(n18), .Z(n729) );
  CNR2XL U880 ( .A(n48), .B(n17), .Z(n742) );
  CNR2XL U881 ( .A(n50), .B(n16), .Z(n756) );
  CNR2XL U882 ( .A(n46), .B(n23), .Z(n674) );
  CNR2XL U883 ( .A(n50), .B(n21), .Z(n691) );
  CNR2XL U884 ( .A(n40), .B(n26), .Z(n656) );
  CNR2XL U885 ( .A(n54), .B(n19), .Z(n712) );
  CNR2XL U886 ( .A(n34), .B(n15), .Z(n779) );
  CNR2XL U887 ( .A(n40), .B(n54), .Z(n826) );
  CNR2XL U888 ( .A(n54), .B(n16), .Z(n754) );
  CNR2XL U889 ( .A(n42), .B(n22), .Z(n685) );
  CNR2XL U890 ( .A(n38), .B(n22), .Z(n687) );
  CNR2XL U891 ( .A(n44), .B(n19), .Z(n717) );
  CNR2XL U892 ( .A(n46), .B(n21), .Z(n693) );
  CEOXL U893 ( .A(n213), .B(n1000), .Z(product[3]) );
  CNR2XL U894 ( .A(n38), .B(n17), .Z(n747) );
  CNR2XL U895 ( .A(n40), .B(n17), .Z(n746) );
  CNR2XL U896 ( .A(n44), .B(n54), .Z(n824) );
  CNR2XL U897 ( .A(n48), .B(n21), .Z(n692) );
  CNR2XL U898 ( .A(n52), .B(n19), .Z(n713) );
  CNR2XL U899 ( .A(n38), .B(n54), .Z(n827) );
  CNR2XL U900 ( .A(n36), .B(n22), .Z(n688) );
  CNR2XL U901 ( .A(n38), .B(n21), .Z(n697) );
  CNR2XL U902 ( .A(n48), .B(n16), .Z(n757) );
  CNR2XL U903 ( .A(n54), .B(n912), .Z(n808) );
  CNR2XL U904 ( .A(n42), .B(n20), .Z(n706) );
  CNR2XL U905 ( .A(n54), .B(n910), .Z(n783) );
  CNR2XL U906 ( .A(n46), .B(n19), .Z(n716) );
  CNR2XL U907 ( .A(n44), .B(n21), .Z(n694) );
  CNR2XL U908 ( .A(n50), .B(n18), .Z(n727) );
  CNR2XL U909 ( .A(n50), .B(n54), .Z(n821) );
  CNR2XL U910 ( .A(n34), .B(n25), .Z(n665) );
  CNR2XL U911 ( .A(n46), .B(n54), .Z(n823) );
  CNR2XL U912 ( .A(n38), .B(n26), .Z(n657) );
  CNR2XL U913 ( .A(n46), .B(n22), .Z(n683) );
  CNR2XL U914 ( .A(n54), .B(n18), .Z(n725) );
  CNR2XL U915 ( .A(n34), .B(n48), .Z(n856) );
  CNR2XL U916 ( .A(n34), .B(n911), .Z(n806) );
  CNR2XL U917 ( .A(n42), .B(n18), .Z(n731) );
  CNR2XL U918 ( .A(n40), .B(n19), .Z(n719) );
  CNR2XL U919 ( .A(n34), .B(n912), .Z(n818) );
  CNR2XL U920 ( .A(n36), .B(n54), .Z(n828) );
  CNR2XL U921 ( .A(n42), .B(n19), .Z(n718) );
  CNR2XL U922 ( .A(n52), .B(n17), .Z(n740) );
  CNR2XL U923 ( .A(n34), .B(n26), .Z(n659) );
  CNR2XL U924 ( .A(n34), .B(n22), .Z(n689) );
  CNR2XL U925 ( .A(n46), .B(n16), .Z(n758) );
  CNR2XL U926 ( .A(n34), .B(n50), .Z(n848) );
  CNR2XL U927 ( .A(n911), .B(n17), .Z(n737) );
  CNR2XL U928 ( .A(n44), .B(n24), .Z(n667) );
  CNR2XL U929 ( .A(n52), .B(n20), .Z(n701) );
  CNR2XL U930 ( .A(n32), .B(n34), .Z(n885) );
  CNR2XL U931 ( .A(n48), .B(n19), .Z(n715) );
  CNR2XL U932 ( .A(n34), .B(n54), .Z(n829) );
  CNR2XL U933 ( .A(n34), .B(n38), .Z(n881) );
  CNR2XL U934 ( .A(n36), .B(n20), .Z(n709) );
  CNR2XL U935 ( .A(n38), .B(n25), .Z(n663) );
  CNR2XL U936 ( .A(n34), .B(n46), .Z(n863) );
  CNR2XL U937 ( .A(n34), .B(n16), .Z(n764) );
  CNR2XL U938 ( .A(n46), .B(n17), .Z(n743) );
  CNR2XL U939 ( .A(n32), .B(n54), .Z(n830) );
  CNR2XL U940 ( .A(n36), .B(n21), .Z(n698) );
  CNR2XL U941 ( .A(n44), .B(n18), .Z(n730) );
  CNR2XL U942 ( .A(n34), .B(n910), .Z(n793) );
  CNR2XL U943 ( .A(n50), .B(n17), .Z(n741) );
  CNR2XL U944 ( .A(n48), .B(n18), .Z(n728) );
  CNR2XL U945 ( .A(n34), .B(n42), .Z(n874) );
  CNR2XL U946 ( .A(n32), .B(n18), .Z(n736) );
  CNR2XL U947 ( .A(n34), .B(n29), .Z(n647) );
  CNR2XL U948 ( .A(n912), .B(n18), .Z(n724) );
  CEO3X1 U949 ( .A(n724), .B(n280), .C(n278), .Z(n248) );
  CNR2XL U950 ( .A(n34), .B(n28), .Z(n650) );
  CNR2XL U951 ( .A(n911), .B(n16), .Z(n752) );
  CNR2XL U952 ( .A(n910), .B(n16), .Z(n751) );
  CEO3X1 U953 ( .A(n661), .B(n652), .C(n656), .Z(n251) );
  CNR2XL U954 ( .A(n48), .B(n22), .Z(n682) );
  CEO3X1 U955 ( .A(n737), .B(n691), .C(n712), .Z(n249) );
  CNR2XL U956 ( .A(n34), .B(n40), .Z(n878) );
  CIVX4 U957 ( .A(b[3]), .Z(n38) );
  CIVX4 U958 ( .A(b[4]), .Z(n40) );
  CNR2XL U959 ( .A(n132), .B(n1041), .Z(n127) );
  CIVX4 U960 ( .A(b[6]), .Z(n44) );
  CIVX4 U961 ( .A(b[5]), .Z(n42) );
  CIVX4 U962 ( .A(b[7]), .Z(n46) );
  CIVX4 U963 ( .A(b[8]), .Z(n48) );
  CIVX3 U964 ( .A(b[12]), .Z(n912) );
  CENX1 U965 ( .A(n991), .B(n85), .Z(product[31]) );
  CENX1 U966 ( .A(n1026), .B(n254), .Z(n991) );
  CND2XL U967 ( .A(n220), .B(n1045), .Z(n65) );
  CNR2XL U968 ( .A(n40), .B(n42), .Z(n871) );
  CIVX1 U969 ( .A(b[28]), .Z(n28) );
  CIVXL U970 ( .A(n1039), .Z(n135) );
  CND2IXL U971 ( .B(n212), .A(n213), .Z(n84) );
  CENX1 U972 ( .A(n77), .B(n186), .Z(product[10]) );
  COND1XL U973 ( .A(n181), .B(n169), .C(n170), .Z(n168) );
  CND2X1 U974 ( .A(n996), .B(n995), .Z(n169) );
  CANR1XL U975 ( .A(n177), .B(n996), .C(n172), .Z(n170) );
  COND1XL U976 ( .A(n166), .B(n162), .C(n163), .Z(n161) );
  COR2X1 U977 ( .A(n549), .B(n562), .Z(n992) );
  CND2XL U978 ( .A(n427), .B(n446), .Z(n108) );
  CND2XL U979 ( .A(n467), .B(n484), .Z(n119) );
  CND2XL U980 ( .A(n447), .B(n466), .Z(n111) );
  COR2X1 U981 ( .A(n519), .B(n534), .Z(n993) );
  COR2X1 U982 ( .A(n485), .B(n502), .Z(n994) );
  CANR1XL U983 ( .A(n194), .B(n999), .C(n191), .Z(n189) );
  COND1XL U984 ( .A(n195), .B(n197), .C(n196), .Z(n194) );
  COND1XL U985 ( .A(n187), .B(n189), .C(n188), .Z(n186) );
  CNR2X1 U986 ( .A(n575), .B(n586), .Z(n162) );
  CENX1 U987 ( .A(n79), .B(n194), .Z(product[8]) );
  CNR2X1 U988 ( .A(n587), .B(n596), .Z(n165) );
  CEOXL U989 ( .A(n189), .B(n78), .Z(product[9]) );
  COR2X1 U990 ( .A(n607), .B(n614), .Z(n995) );
  COR2X1 U991 ( .A(n597), .B(n606), .Z(n996) );
  CND2X1 U992 ( .A(n597), .B(n606), .Z(n174) );
  CND2X1 U993 ( .A(n615), .B(n622), .Z(n185) );
  CND2X1 U994 ( .A(n607), .B(n614), .Z(n179) );
  COR2X1 U995 ( .A(n615), .B(n622), .Z(n997) );
  CND2X1 U996 ( .A(n587), .B(n596), .Z(n166) );
  COR2X1 U997 ( .A(n563), .B(n574), .Z(n998) );
  COND1XL U998 ( .A(n203), .B(n205), .C(n204), .Z(n202) );
  CENX1 U999 ( .A(n81), .B(n202), .Z(product[6]) );
  CENX1 U1000 ( .A(n93), .B(n60), .Z(product[27]) );
  CND2X1 U1001 ( .A(n1003), .B(n92), .Z(n60) );
  CNR2X1 U1002 ( .A(n635), .B(n638), .Z(n195) );
  CNR2X1 U1003 ( .A(n623), .B(n628), .Z(n187) );
  CEOXL U1004 ( .A(n205), .B(n82), .Z(product[5]) );
  CND2X1 U1005 ( .A(n629), .B(n634), .Z(n193) );
  CND2X1 U1006 ( .A(n635), .B(n638), .Z(n196) );
  CND2X1 U1007 ( .A(n623), .B(n628), .Z(n188) );
  COR2X1 U1008 ( .A(n629), .B(n634), .Z(n999) );
  CENX1 U1009 ( .A(n83), .B(n210), .Z(product[4]) );
  CNR2X1 U1010 ( .A(n213), .B(n1000), .Z(n210) );
  CNR2X1 U1011 ( .A(n40), .B(n46), .Z(n860) );
  CNR2X1 U1012 ( .A(n42), .B(n24), .Z(n668) );
  CNR2X1 U1013 ( .A(n40), .B(n48), .Z(n853) );
  CNR2X1 U1014 ( .A(n48), .B(n911), .Z(n799) );
  CNR2X1 U1015 ( .A(n50), .B(n912), .Z(n810) );
  CNR2X1 U1016 ( .A(n54), .B(n52), .Z(n820) );
  CNR2X1 U1017 ( .A(n38), .B(n911), .Z(n804) );
  CNR2X1 U1018 ( .A(n32), .B(n16), .Z(n765) );
  CNR2X1 U1019 ( .A(n54), .B(n42), .Z(n825) );
  CNR2X1 U1020 ( .A(n911), .B(n910), .Z(n781) );
  CNR2X1 U1021 ( .A(n40), .B(n23), .Z(n677) );
  CENX1 U1022 ( .A(n101), .B(n62), .Z(product[25]) );
  CND2X1 U1023 ( .A(n1005), .B(n100), .Z(n62) );
  CNR2X1 U1024 ( .A(n911), .B(n42), .Z(n802) );
  CNR2X1 U1025 ( .A(n48), .B(n50), .Z(n841) );
  CNR2X1 U1026 ( .A(n40), .B(n911), .Z(n803) );
  CNR2X1 U1027 ( .A(n912), .B(n42), .Z(n814) );
  CNR2X1 U1028 ( .A(n46), .B(n910), .Z(n787) );
  CNR2X1 U1029 ( .A(n44), .B(n15), .Z(n774) );
  CNR2X1 U1030 ( .A(n38), .B(n18), .Z(n733) );
  CNR2X1 U1031 ( .A(n42), .B(n23), .Z(n676) );
  CNR2X1 U1032 ( .A(n46), .B(n48), .Z(n850) );
  CNR2X1 U1033 ( .A(n52), .B(n15), .Z(n770) );
  CNR2X1 U1034 ( .A(n44), .B(n48), .Z(n851) );
  CNR2X1 U1035 ( .A(n643), .B(n644), .Z(n203) );
  CNR2X1 U1036 ( .A(n50), .B(n910), .Z(n785) );
  CNR2X1 U1037 ( .A(n36), .B(n19), .Z(n721) );
  CNR2X1 U1038 ( .A(n42), .B(n16), .Z(n760) );
  CNR2X1 U1039 ( .A(n32), .B(n21), .Z(n700) );
  CNR2X1 U1040 ( .A(n48), .B(n52), .Z(n832) );
  CNR2X1 U1041 ( .A(n44), .B(n911), .Z(n801) );
  CNR2X1 U1042 ( .A(n46), .B(n912), .Z(n812) );
  CNR2X1 U1043 ( .A(n50), .B(n52), .Z(n831) );
  CNR2X1 U1044 ( .A(n46), .B(n50), .Z(n842) );
  CNR2X1 U1045 ( .A(n44), .B(n52), .Z(n834) );
  CNR2X1 U1046 ( .A(n38), .B(n910), .Z(n791) );
  CNR2X1 U1047 ( .A(n40), .B(n24), .Z(n669) );
  CNR2X1 U1048 ( .A(n44), .B(n46), .Z(n858) );
  CNR2X1 U1049 ( .A(n38), .B(n52), .Z(n837) );
  CNR2X1 U1050 ( .A(n912), .B(n911), .Z(n795) );
  CNR2X1 U1051 ( .A(n52), .B(n16), .Z(n755) );
  CNR2X1 U1052 ( .A(n42), .B(n21), .Z(n695) );
  CNR2X1 U1053 ( .A(n48), .B(n910), .Z(n786) );
  CNR2X1 U1054 ( .A(n912), .B(n52), .Z(n809) );
  CNR2X1 U1055 ( .A(n40), .B(n18), .Z(n732) );
  CNR2X1 U1056 ( .A(n40), .B(n44), .Z(n866) );
  CNR2X1 U1057 ( .A(n38), .B(n46), .Z(n861) );
  CNR2X1 U1058 ( .A(n38), .B(n48), .Z(n854) );
  CNR2X1 U1059 ( .A(n911), .B(n15), .Z(n767) );
  CNR2X1 U1060 ( .A(n48), .B(n20), .Z(n703) );
  CNR2X1 U1061 ( .A(n34), .B(n27), .Z(n654) );
  CNR2X1 U1062 ( .A(n38), .B(n19), .Z(n720) );
  CNR2X1 U1063 ( .A(n32), .B(n22), .Z(n690) );
  CNR2X1 U1064 ( .A(n34), .B(n21), .Z(n699) );
  CNR2X1 U1065 ( .A(n38), .B(n42), .Z(n872) );
  CNR2X1 U1066 ( .A(n50), .B(n42), .Z(n844) );
  CEOXL U1067 ( .A(n61), .B(n96), .Z(product[26]) );
  CND2X1 U1068 ( .A(n216), .B(n95), .Z(n61) );
  CNR2X1 U1069 ( .A(n912), .B(n16), .Z(n753) );
  CNR2X1 U1070 ( .A(n44), .B(n22), .Z(n684) );
  CNR2X1 U1071 ( .A(n32), .B(n23), .Z(n681) );
  CNR2X1 U1072 ( .A(n48), .B(n912), .Z(n811) );
  CNR2X1 U1073 ( .A(n36), .B(n18), .Z(n734) );
  CNR2X1 U1074 ( .A(n34), .B(n19), .Z(n722) );
  CNR2X1 U1075 ( .A(n32), .B(n24), .Z(n673) );
  CNR2X1 U1076 ( .A(n44), .B(n50), .Z(n843) );
  CNR2X1 U1077 ( .A(n40), .B(n15), .Z(n776) );
  CNR2X1 U1078 ( .A(n36), .B(n17), .Z(n748) );
  CNR2X1 U1079 ( .A(n910), .B(n42), .Z(n789) );
  COR2X1 U1080 ( .A(n645), .B(n882), .Z(n1001) );
  CNR2X1 U1081 ( .A(n50), .B(n911), .Z(n798) );
  CAOR1X1 U1082 ( .A(n1003), .B(n93), .C(n90), .Z(n1002) );
  CNR2X1 U1083 ( .A(n38), .B(n24), .Z(n670) );
  CNR2X1 U1084 ( .A(n44), .B(n912), .Z(n813) );
  CNR2X1 U1085 ( .A(n38), .B(n15), .Z(n777) );
  CNR2X1 U1086 ( .A(n40), .B(n50), .Z(n845) );
  CNR2X1 U1087 ( .A(n38), .B(n23), .Z(n678) );
  CNR2X1 U1088 ( .A(n32), .B(n19), .Z(n723) );
  CNR2X1 U1089 ( .A(n38), .B(n16), .Z(n762) );
  CNR2X1 U1090 ( .A(n38), .B(n50), .Z(n846) );
  CNR2X1 U1091 ( .A(n32), .B(n46), .Z(n864) );
  CNR2X1 U1092 ( .A(n48), .B(n15), .Z(n772) );
  CNR2X1 U1093 ( .A(n911), .B(n52), .Z(n797) );
  CNR2X1 U1094 ( .A(n54), .B(n15), .Z(n769) );
  CNR2X1 U1095 ( .A(n32), .B(n26), .Z(n660) );
  CNR2X1 U1096 ( .A(n44), .B(n20), .Z(n705) );
  CNR2X1 U1097 ( .A(n46), .B(n911), .Z(n800) );
  CNR2X1 U1098 ( .A(n44), .B(n910), .Z(n788) );
  CNR2X1 U1099 ( .A(n40), .B(n16), .Z(n761) );
  CNR2X1 U1100 ( .A(n910), .B(n15), .Z(n766) );
  CNR2X1 U1101 ( .A(n50), .B(n20), .Z(n702) );
  CNR2X1 U1102 ( .A(n32), .B(n29), .Z(n648) );
  CNR2X1 U1103 ( .A(n50), .B(n15), .Z(n771) );
  CNR2X1 U1104 ( .A(n910), .B(n52), .Z(n784) );
  CNR2X1 U1105 ( .A(n44), .B(n16), .Z(n759) );
  CNR2X1 U1106 ( .A(n46), .B(n15), .Z(n773) );
  CNR2X1 U1107 ( .A(n54), .B(n911), .Z(n796) );
  CNR2X1 U1108 ( .A(n40), .B(n20), .Z(n707) );
  CEOX1 U1109 ( .A(n646), .B(n647), .Z(n253) );
  CND2X1 U1110 ( .A(n645), .B(n882), .Z(n209) );
  CND2X1 U1111 ( .A(n639), .B(n641), .Z(n201) );
  CND2X1 U1112 ( .A(n335), .B(n358), .Z(n92) );
  CNR2X1 U1113 ( .A(n44), .B(n23), .Z(n675) );
  CND2X1 U1114 ( .A(n643), .B(n644), .Z(n204) );
  COR2X1 U1115 ( .A(n335), .B(n358), .Z(n1003) );
  COR2X1 U1116 ( .A(n639), .B(n641), .Z(n1004) );
  CEOXL U1117 ( .A(n63), .B(n104), .Z(product[24]) );
  CND2X1 U1118 ( .A(n218), .B(n103), .Z(n63) );
  CNR2XL U1119 ( .A(n1048), .B(n1046), .Z(n105) );
  COND1XL U1120 ( .A(n1045), .B(n1048), .C(n1047), .Z(n106) );
  CIVX4 U1121 ( .A(b[1]), .Z(n34) );
  CND2XL U1122 ( .A(n1053), .B(n1052), .Z(n147) );
  CANR1XL U1123 ( .A(n155), .B(n1053), .C(n150), .Z(n148) );
  CND2XL U1124 ( .A(n221), .B(n1055), .Z(n114) );
  CANR1XL U1125 ( .A(n122), .B(n221), .C(n117), .Z(n115) );
  CANR1XL U1126 ( .A(n142), .B(n1054), .C(n135), .Z(n133) );
  CIVX2 U1127 ( .A(b[21]), .Z(n21) );
  CIVX2 U1128 ( .A(b[11]), .Z(n54) );
  CIVX2 U1129 ( .A(b[22]), .Z(n22) );
  CIVX2 U1130 ( .A(b[16]), .Z(n16) );
  CENX1 U1131 ( .A(n109), .B(n64), .Z(product[23]) );
  CND2XL U1132 ( .A(n219), .B(n1047), .Z(n64) );
  COND1XL U1133 ( .A(n1046), .B(n112), .C(n1045), .Z(n109) );
  CNR2X1 U1134 ( .A(n1007), .B(n1006), .Z(n102) );
  CNR2X1 U1135 ( .A(n359), .B(n1011), .Z(n94) );
  CIVX2 U1136 ( .A(b[18]), .Z(n18) );
  CNR2XL U1137 ( .A(n38), .B(n20), .Z(n708) );
  CNR2XL U1138 ( .A(n32), .B(n42), .Z(n875) );
  CNR2XL U1139 ( .A(n34), .B(n52), .Z(n839) );
  CIVX2 U1140 ( .A(b[19]), .Z(n19) );
  CIVX2 U1141 ( .A(b[20]), .Z(n20) );
  COR2X1 U1142 ( .A(n1010), .B(n1008), .Z(n1005) );
  CNR2X1 U1143 ( .A(n34), .B(n20), .Z(n710) );
  CNR2XL U1144 ( .A(n40), .B(n25), .Z(n662) );
  CNR2X1 U1145 ( .A(n46), .B(n20), .Z(n704) );
  CNR2XL U1146 ( .A(n34), .B(n18), .Z(n735) );
  CNR2XL U1147 ( .A(n48), .B(n42), .Z(n852) );
  CNR2XL U1148 ( .A(n32), .B(n25), .Z(n666) );
  CNR2XL U1149 ( .A(n36), .B(n42), .Z(n873) );
  CNR2XL U1150 ( .A(n32), .B(n15), .Z(n780) );
  CND2X1 U1151 ( .A(n1010), .B(n1008), .Z(n100) );
  CND2X1 U1152 ( .A(n1007), .B(n1006), .Z(n103) );
  CND2X1 U1153 ( .A(n359), .B(n1011), .Z(n95) );
  CEOX1 U1154 ( .A(n66), .B(n120), .Z(product[21]) );
  CND2XL U1155 ( .A(n221), .B(n1043), .Z(n66) );
  CANR1XL U1156 ( .A(n1055), .B(n125), .C(n122), .Z(n120) );
  CEOX1 U1157 ( .A(n71), .B(n153), .Z(product[16]) );
  CND2XL U1158 ( .A(n1053), .B(n1036), .Z(n71) );
  CANR1XL U1159 ( .A(n1052), .B(n158), .C(n155), .Z(n153) );
  CENX1 U1160 ( .A(n131), .B(n68), .Z(product[19]) );
  CND2XL U1161 ( .A(n223), .B(n1040), .Z(n68) );
  COND1XL U1162 ( .A(n132), .B(n145), .C(n133), .Z(n131) );
  CENX1 U1163 ( .A(n138), .B(n69), .Z(product[18]) );
  CND2XL U1164 ( .A(n1054), .B(n1039), .Z(n69) );
  COND1XL U1165 ( .A(n1038), .B(n145), .C(n1037), .Z(n138) );
  CENX1 U1166 ( .A(n164), .B(n1033), .Z(n1087) );
  COND1XL U1167 ( .A(n1032), .B(n167), .C(n1031), .Z(n164) );
  CENX1 U1168 ( .A(n125), .B(n67), .Z(product[20]) );
  CND2XL U1169 ( .A(n1055), .B(n1042), .Z(n67) );
  CENX1 U1170 ( .A(n158), .B(n72), .Z(product[15]) );
  CND2XL U1171 ( .A(n1052), .B(n1035), .Z(n72) );
  CENX1 U1172 ( .A(n1029), .B(n1049), .Z(n1089) );
  CEOX1 U1173 ( .A(n175), .B(n1030), .Z(n1088) );
  CANR1XL U1174 ( .A(n1051), .B(n1049), .C(n1050), .Z(n175) );
  CEOX1 U1175 ( .A(n65), .B(n112), .Z(product[22]) );
  CEOX1 U1176 ( .A(n70), .B(n145), .Z(product[17]) );
  CND2XL U1177 ( .A(n225), .B(n1037), .Z(n70) );
  CEOX1 U1178 ( .A(n74), .B(n167), .Z(product[13]) );
  CND2X1 U1179 ( .A(n229), .B(n1031), .Z(n74) );
  CNR2XL U1180 ( .A(n885), .B(a[1]), .Z(n212) );
  CIVX2 U1181 ( .A(n84), .Z(product[2]) );
  CIVX2 U1182 ( .A(n100), .Z(n98) );
  CIVX2 U1183 ( .A(n92), .Z(n90) );
  CIVX2 U1184 ( .A(b[30]), .Z(n30) );
  CIVX2 U1185 ( .A(b[29]), .Z(n29) );
  CIVX2 U1186 ( .A(b[27]), .Z(n27) );
  CIVX2 U1187 ( .A(b[26]), .Z(n26) );
  CIVX2 U1188 ( .A(b[25]), .Z(n25) );
  CIVX2 U1189 ( .A(n203), .Z(n237) );
  CIVX2 U1190 ( .A(n195), .Z(n235) );
  CIVX2 U1191 ( .A(n187), .Z(n233) );
  CIVX2 U1192 ( .A(b[23]), .Z(n23) );
  CIVX2 U1193 ( .A(n1032), .Z(n229) );
  CIVX2 U1194 ( .A(n1041), .Z(n223) );
  CIVX2 U1195 ( .A(n1046), .Z(n220) );
  CIVX2 U1196 ( .A(n1048), .Z(n219) );
  CIVX2 U1197 ( .A(n102), .Z(n218) );
  CIVX2 U1198 ( .A(n94), .Z(n216) );
  CIVX2 U1199 ( .A(n209), .Z(n207) );
  CIVX2 U1200 ( .A(n201), .Z(n199) );
  CIVX2 U1201 ( .A(n193), .Z(n191) );
  CIVX2 U1202 ( .A(n185), .Z(n183) );
  CIVX2 U1203 ( .A(n174), .Z(n172) );
  CIVX2 U1204 ( .A(n1027), .Z(n167) );
  CIVX2 U1205 ( .A(n159), .Z(n158) );
  CIVX2 U1206 ( .A(n1035), .Z(n155) );
  CIVX2 U1207 ( .A(n146), .Z(n145) );
  CIVX2 U1208 ( .A(n1037), .Z(n142) );
  CIVX2 U1209 ( .A(n1038), .Z(n225) );
  CIVX2 U1210 ( .A(n1042), .Z(n122) );
  CIVX2 U1211 ( .A(n1043), .Z(n117) );
  CIVX2 U1212 ( .A(n1044), .Z(n221) );
  CIVX2 U1213 ( .A(n113), .Z(n112) );
endmodule


module calc_DW02_mult_2_stage_10 ( A, B, TC, CLK, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC, CLK;
  wire   n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, \B_extended[32] ,
         n6, n8, n10, n12, n14, n16, n18, n20, n22, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34;
  assign \B_extended[32]  = B[31];

  calc_DW_mult_tc_21 mult_96 ( .a({\B_extended[32] , A}), .b({\B_extended[32] , 
        \B_extended[32] , B[30:0]}), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, PRODUCT[31:11], n35, n36, n37, n38, n39, n40, 
        n41, n42, n43, SYNOPSYS_UNCONNECTED__34, n44}), .dw1_CLK(CLK) );
  CFD1QXL clk_r_REG56_S1 ( .D(n43), .CP(CLK), .Q(n26) );
  CFD1QXL clk_r_REG57_S1 ( .D(n42), .CP(CLK), .Q(n27) );
  CFD1QXL clk_r_REG55_S1 ( .D(n40), .CP(CLK), .Q(n29) );
  CFD1QXL clk_r_REG52_S1 ( .D(n39), .CP(CLK), .Q(n30) );
  CFD1QXL clk_r_REG54_S1 ( .D(n41), .CP(CLK), .Q(n28) );
  CFD1QXL clk_r_REG51_S1 ( .D(n36), .CP(CLK), .Q(n33) );
  CFD1QXL clk_r_REG53_S1 ( .D(n38), .CP(CLK), .Q(n31) );
  CFD1QXL clk_r_REG50_S1 ( .D(n37), .CP(CLK), .Q(n32) );
  CFD1QXL clk_r_REG45_S1 ( .D(n35), .CP(CLK), .Q(n34) );
  CFD1QXL clk_r_REG59_S1 ( .D(n44), .CP(CLK), .Q(n25) );
  CIVDX1 U1 ( .A(n29), .Z1(n8) );
  CIVDXL U2 ( .A(n31), .Z1(n6) );
  CNIVX1 U3 ( .A(n6), .Z(PRODUCT[7]) );
  CNIVX1 U4 ( .A(n8), .Z(PRODUCT[5]) );
  CIVDXL U5 ( .A(n27), .Z1(n10) );
  CNIVX1 U6 ( .A(n10), .Z(PRODUCT[3]) );
  CIVDXL U7 ( .A(n33), .Z1(n12) );
  CNIVX1 U8 ( .A(n12), .Z(PRODUCT[9]) );
  CIVDX1 U9 ( .A(n26), .Z1(n14) );
  CNIVX1 U10 ( .A(n14), .Z(PRODUCT[2]) );
  CIVDX1 U11 ( .A(n25), .Z1(n16) );
  CNIVX1 U12 ( .A(n16), .Z(PRODUCT[0]) );
  CIVDX1 U13 ( .A(n28), .Z1(n18) );
  CNIVX1 U14 ( .A(n18), .Z(PRODUCT[4]) );
  CIVDX1 U15 ( .A(n30), .Z1(n20) );
  CNIVX1 U16 ( .A(n20), .Z(PRODUCT[6]) );
  CIVDX1 U17 ( .A(n32), .Z1(n22) );
  CNIVX1 U18 ( .A(n22), .Z(PRODUCT[8]) );
  CIVDX1 U19 ( .A(n34), .Z1(n24) );
  CNIVX1 U20 ( .A(n24), .Z(PRODUCT[10]) );
endmodule


module calc_DW01_add_6 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n38, n40, n41, n42, n43, n44, n46, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n62, n64,
         n65, n66, n67, n68, n69, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n204, n206, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n335, n336, n337, n338;

  CANR1X1 U268 ( .A(n338), .B(n41), .C(n38), .Z(n36) );
  CENXL U269 ( .A(n41), .B(n3), .Z(SUM[29]) );
  COND1X1 U270 ( .A(n42), .B(n44), .C(n43), .Z(n41) );
  COND1X1 U271 ( .A(n50), .B(n117), .C(n51), .Z(n49) );
  CIVX1 U272 ( .A(n117), .Z(n116) );
  CANR1X1 U273 ( .A(n167), .B(n118), .C(n119), .Z(n117) );
  CNR2XL U274 ( .A(n141), .B(n136), .Z(n134) );
  CNR2XL U275 ( .A(A[12]), .B(B[12]), .Z(n141) );
  CND2XL U276 ( .A(A[2]), .B(B[2]), .Z(n195) );
  CNR2XL U277 ( .A(n154), .B(n149), .Z(n147) );
  CNR2XL U278 ( .A(n129), .B(n124), .Z(n122) );
  CND2XL U279 ( .A(A[23]), .B(B[23]), .Z(n81) );
  CND2XL U280 ( .A(A[21]), .B(B[21]), .Z(n89) );
  CANR1XL U281 ( .A(n95), .B(n116), .C(n96), .Z(n94) );
  CND2X1 U282 ( .A(n86), .B(n78), .Z(n76) );
  CNR2X1 U283 ( .A(n114), .B(n109), .Z(n107) );
  CNR2X1 U284 ( .A(n185), .B(n180), .Z(n178) );
  CANR1XL U285 ( .A(n197), .B(n189), .C(n190), .Z(n188) );
  CNR2X1 U286 ( .A(n91), .B(n88), .Z(n86) );
  CNR2X1 U287 ( .A(A[16]), .B(B[16]), .Z(n114) );
  CIVXL U288 ( .A(n73), .Z(n72) );
  CIVXL U289 ( .A(n144), .Z(n143) );
  CIVXL U290 ( .A(n98), .Z(n96) );
  CNR2XL U291 ( .A(n194), .B(n191), .Z(n189) );
  CIVXL U292 ( .A(n64), .Z(n62) );
  CNR2XL U293 ( .A(n164), .B(n161), .Z(n159) );
  CNR2XL U294 ( .A(n104), .B(n101), .Z(n99) );
  CND2XL U295 ( .A(n68), .B(n336), .Z(n59) );
  CIVXL U296 ( .A(n185), .Z(n228) );
  CIVX1 U297 ( .A(n54), .Z(n206) );
  CND2XL U298 ( .A(n229), .B(n192), .Z(n29) );
  CNR2XL U299 ( .A(A[8]), .B(B[8]), .Z(n164) );
  CNR2XL U300 ( .A(A[24]), .B(B[24]), .Z(n66) );
  CND2XL U301 ( .A(A[6]), .B(B[6]), .Z(n176) );
  CND2XL U302 ( .A(A[18]), .B(B[18]), .Z(n105) );
  CND2XL U303 ( .A(A[1]), .B(B[1]), .Z(n199) );
  CND2XL U304 ( .A(A[26]), .B(B[26]), .Z(n55) );
  CENX1 U305 ( .A(n335), .B(n33), .Z(SUM[31]) );
  CENX1 U306 ( .A(B[31]), .B(A[31]), .Z(n335) );
  CND2XL U307 ( .A(n209), .B(n81), .Z(n9) );
  CEOXL U308 ( .A(n2), .B(n36), .Z(SUM[30]) );
  CEOXL U309 ( .A(n17), .B(n126), .Z(SUM[15]) );
  CND2XL U310 ( .A(n217), .B(n125), .Z(n17) );
  CND2XL U311 ( .A(n210), .B(n84), .Z(n10) );
  CEOXL U312 ( .A(n10), .B(n85), .Z(SUM[22]) );
  CEOXL U313 ( .A(n6), .B(n56), .Z(SUM[26]) );
  CEOXL U314 ( .A(n4), .B(n44), .Z(SUM[28]) );
  CND2XL U315 ( .A(n336), .B(n64), .Z(n7) );
  CND2XL U316 ( .A(n68), .B(n67), .Z(n8) );
  CND2XL U317 ( .A(n211), .B(n89), .Z(n11) );
  CND2XL U318 ( .A(n212), .B(n92), .Z(n12) );
  CND2XL U319 ( .A(n213), .B(n102), .Z(n13) );
  CND2XL U320 ( .A(n214), .B(n105), .Z(n14) );
  CND2XL U321 ( .A(n215), .B(n110), .Z(n15) );
  CND2XL U322 ( .A(n216), .B(n115), .Z(n16) );
  CND2XL U323 ( .A(n218), .B(n130), .Z(n18) );
  CND2XL U324 ( .A(n219), .B(n137), .Z(n19) );
  CND2XL U325 ( .A(n220), .B(n142), .Z(n20) );
  CEOXL U326 ( .A(n20), .B(n143), .Z(SUM[12]) );
  CND2XL U327 ( .A(n221), .B(n150), .Z(n21) );
  CND2XL U328 ( .A(n222), .B(n155), .Z(n22) );
  CND2XL U329 ( .A(n223), .B(n162), .Z(n23) );
  CND2XL U330 ( .A(n224), .B(n165), .Z(n24) );
  CEOXL U331 ( .A(n24), .B(n166), .Z(SUM[8]) );
  CND2XL U332 ( .A(n225), .B(n173), .Z(n25) );
  CND2XL U333 ( .A(n226), .B(n176), .Z(n26) );
  CND2XL U334 ( .A(n227), .B(n181), .Z(n27) );
  CND2XL U335 ( .A(n228), .B(n186), .Z(n28) );
  CND2XL U336 ( .A(n230), .B(n195), .Z(n30) );
  CND2XL U337 ( .A(n231), .B(n199), .Z(n31) );
  CEOXL U338 ( .A(n201), .B(n31), .Z(SUM[1]) );
  CND2IXL U339 ( .B(n200), .A(n201), .Z(n32) );
  CNR2X1 U340 ( .A(n97), .B(n76), .Z(n74) );
  CANR1XL U341 ( .A(n86), .B(n93), .C(n87), .Z(n85) );
  CANR1XL U342 ( .A(n107), .B(n116), .C(n108), .Z(n106) );
  CANR1XL U343 ( .A(n178), .B(n187), .C(n179), .Z(n177) );
  COND1XL U344 ( .A(n132), .B(n143), .C(n133), .Z(n131) );
  COND1XL U345 ( .A(n157), .B(n166), .C(n158), .Z(n156) );
  CNR2X1 U346 ( .A(n145), .B(n120), .Z(n118) );
  COND1XL U347 ( .A(n120), .B(n146), .C(n121), .Z(n119) );
  CND2X1 U348 ( .A(n134), .B(n122), .Z(n120) );
  CANR1XL U349 ( .A(n74), .B(n116), .C(n75), .Z(n73) );
  COND1XL U350 ( .A(n145), .B(n166), .C(n146), .Z(n144) );
  CND2X1 U351 ( .A(n107), .B(n99), .Z(n97) );
  CND2X1 U352 ( .A(n159), .B(n147), .Z(n145) );
  CANR1XL U353 ( .A(n337), .B(n49), .C(n46), .Z(n44) );
  CND2X1 U354 ( .A(n74), .B(n52), .Z(n50) );
  CANR1XL U355 ( .A(n52), .B(n75), .C(n53), .Z(n51) );
  CNR2X1 U356 ( .A(n59), .B(n54), .Z(n52) );
  CANR1XL U357 ( .A(n69), .B(n336), .C(n62), .Z(n60) );
  COND1XL U358 ( .A(n195), .B(n191), .C(n192), .Z(n190) );
  CANR1XL U359 ( .A(n108), .B(n99), .C(n100), .Z(n98) );
  COND1XL U360 ( .A(n105), .B(n101), .C(n102), .Z(n100) );
  COND1XL U361 ( .A(n201), .B(n198), .C(n199), .Z(n197) );
  COND1XL U362 ( .A(n165), .B(n161), .C(n162), .Z(n160) );
  COND1XL U363 ( .A(n142), .B(n136), .C(n137), .Z(n135) );
  COND1XL U364 ( .A(n168), .B(n188), .C(n169), .Z(n167) );
  CND2X1 U365 ( .A(n178), .B(n170), .Z(n168) );
  CANR1XL U366 ( .A(n179), .B(n170), .C(n171), .Z(n169) );
  CNR2X1 U367 ( .A(n175), .B(n172), .Z(n170) );
  CANR1XL U368 ( .A(n160), .B(n147), .C(n148), .Z(n146) );
  COND1XL U369 ( .A(n155), .B(n149), .C(n150), .Z(n148) );
  COND1XL U370 ( .A(n186), .B(n180), .C(n181), .Z(n179) );
  COND1XL U371 ( .A(n115), .B(n109), .C(n110), .Z(n108) );
  COND1XL U372 ( .A(n92), .B(n88), .C(n89), .Z(n87) );
  COND1XL U373 ( .A(n76), .B(n98), .C(n77), .Z(n75) );
  CANR1XL U374 ( .A(n87), .B(n78), .C(n79), .Z(n77) );
  COND1XL U375 ( .A(n84), .B(n80), .C(n81), .Z(n79) );
  CANR1XL U376 ( .A(n135), .B(n122), .C(n123), .Z(n121) );
  COND1XL U377 ( .A(n130), .B(n124), .C(n125), .Z(n123) );
  CNR2X1 U378 ( .A(n83), .B(n80), .Z(n78) );
  COND1XL U379 ( .A(n54), .B(n60), .C(n55), .Z(n53) );
  COND1XL U380 ( .A(n176), .B(n172), .C(n173), .Z(n171) );
  CNR2X1 U381 ( .A(A[26]), .B(B[26]), .Z(n54) );
  CNR2X1 U382 ( .A(A[5]), .B(B[5]), .Z(n180) );
  CNR2X1 U383 ( .A(A[7]), .B(B[7]), .Z(n172) );
  CNR2X1 U384 ( .A(A[15]), .B(B[15]), .Z(n124) );
  CNR2X1 U385 ( .A(A[13]), .B(B[13]), .Z(n136) );
  CNR2X1 U386 ( .A(A[11]), .B(B[11]), .Z(n149) );
  CNR2X1 U387 ( .A(A[9]), .B(B[9]), .Z(n161) );
  CNR2X1 U388 ( .A(A[23]), .B(B[23]), .Z(n80) );
  CNR2X1 U389 ( .A(A[21]), .B(B[21]), .Z(n88) );
  CNR2X1 U390 ( .A(A[19]), .B(B[19]), .Z(n101) );
  CNR2X1 U391 ( .A(A[17]), .B(B[17]), .Z(n109) );
  CNR2X1 U392 ( .A(A[3]), .B(B[3]), .Z(n191) );
  CNR2X1 U393 ( .A(A[22]), .B(B[22]), .Z(n83) );
  CNR2X1 U394 ( .A(A[18]), .B(B[18]), .Z(n104) );
  CNR2X1 U395 ( .A(A[6]), .B(B[6]), .Z(n175) );
  CNR2X1 U396 ( .A(A[2]), .B(B[2]), .Z(n194) );
  CNR2X1 U397 ( .A(A[20]), .B(B[20]), .Z(n91) );
  CNR2X1 U398 ( .A(A[14]), .B(B[14]), .Z(n129) );
  CNR2X1 U399 ( .A(A[10]), .B(B[10]), .Z(n154) );
  CNR2X1 U400 ( .A(A[4]), .B(B[4]), .Z(n185) );
  CND2X1 U401 ( .A(A[0]), .B(B[0]), .Z(n201) );
  CNR2X1 U402 ( .A(A[28]), .B(B[28]), .Z(n42) );
  CNR2X1 U403 ( .A(A[1]), .B(B[1]), .Z(n198) );
  COR2X1 U404 ( .A(A[25]), .B(B[25]), .Z(n336) );
  CND2X1 U405 ( .A(A[24]), .B(B[24]), .Z(n67) );
  CND2X1 U406 ( .A(A[4]), .B(B[4]), .Z(n186) );
  CND2X1 U407 ( .A(A[10]), .B(B[10]), .Z(n155) );
  CND2X1 U408 ( .A(A[14]), .B(B[14]), .Z(n130) );
  CND2X1 U409 ( .A(A[12]), .B(B[12]), .Z(n142) );
  CND2X1 U410 ( .A(A[16]), .B(B[16]), .Z(n115) );
  CND2X1 U411 ( .A(A[22]), .B(B[22]), .Z(n84) );
  CND2X1 U412 ( .A(A[20]), .B(B[20]), .Z(n92) );
  CND2X1 U413 ( .A(A[8]), .B(B[8]), .Z(n165) );
  CND2X1 U414 ( .A(A[25]), .B(B[25]), .Z(n64) );
  CND2X1 U415 ( .A(A[27]), .B(B[27]), .Z(n48) );
  CND2XL U416 ( .A(A[19]), .B(B[19]), .Z(n102) );
  CND2XL U417 ( .A(A[17]), .B(B[17]), .Z(n110) );
  CND2XL U418 ( .A(A[15]), .B(B[15]), .Z(n125) );
  CND2XL U419 ( .A(A[13]), .B(B[13]), .Z(n137) );
  CND2XL U420 ( .A(A[11]), .B(B[11]), .Z(n150) );
  CND2XL U421 ( .A(A[9]), .B(B[9]), .Z(n162) );
  CND2XL U422 ( .A(A[7]), .B(B[7]), .Z(n173) );
  CND2XL U423 ( .A(A[5]), .B(B[5]), .Z(n181) );
  CND2XL U424 ( .A(A[3]), .B(B[3]), .Z(n192) );
  CND2X1 U425 ( .A(A[28]), .B(B[28]), .Z(n43) );
  COR2X1 U426 ( .A(A[27]), .B(B[27]), .Z(n337) );
  COND1XL U427 ( .A(n34), .B(n36), .C(n35), .Z(n33) );
  CND2X1 U428 ( .A(n202), .B(n35), .Z(n2) );
  CND2X1 U429 ( .A(n338), .B(n40), .Z(n3) );
  CND2X1 U430 ( .A(n204), .B(n43), .Z(n4) );
  CENX1 U431 ( .A(n49), .B(n5), .Z(SUM[27]) );
  CND2X1 U432 ( .A(n337), .B(n48), .Z(n5) );
  CND2X1 U433 ( .A(n206), .B(n55), .Z(n6) );
  CANR1XL U434 ( .A(n57), .B(n72), .C(n58), .Z(n56) );
  CENX1 U435 ( .A(n65), .B(n7), .Z(SUM[25]) );
  COND1XL U436 ( .A(n66), .B(n73), .C(n67), .Z(n65) );
  CENX1 U437 ( .A(n72), .B(n8), .Z(SUM[24]) );
  CENX1 U438 ( .A(n82), .B(n9), .Z(SUM[23]) );
  COND1XL U439 ( .A(n83), .B(n85), .C(n84), .Z(n82) );
  CENX1 U440 ( .A(n90), .B(n11), .Z(SUM[21]) );
  COND1XL U441 ( .A(n91), .B(n94), .C(n92), .Z(n90) );
  CENX1 U442 ( .A(n93), .B(n12), .Z(SUM[20]) );
  CENX1 U443 ( .A(n103), .B(n13), .Z(SUM[19]) );
  COND1XL U444 ( .A(n104), .B(n106), .C(n105), .Z(n103) );
  CEOX1 U445 ( .A(n14), .B(n106), .Z(SUM[18]) );
  CEOX1 U446 ( .A(n15), .B(n111), .Z(SUM[17]) );
  CANR1XL U447 ( .A(n216), .B(n116), .C(n113), .Z(n111) );
  CENX1 U448 ( .A(n116), .B(n16), .Z(SUM[16]) );
  CANR1XL U449 ( .A(n218), .B(n131), .C(n128), .Z(n126) );
  CENX1 U450 ( .A(n131), .B(n18), .Z(SUM[14]) );
  CEOX1 U451 ( .A(n19), .B(n138), .Z(SUM[13]) );
  CANR1XL U452 ( .A(n220), .B(n144), .C(n140), .Z(n138) );
  CEOX1 U453 ( .A(n21), .B(n151), .Z(SUM[11]) );
  CANR1XL U454 ( .A(n222), .B(n156), .C(n153), .Z(n151) );
  CENX1 U455 ( .A(n156), .B(n22), .Z(SUM[10]) );
  CENX1 U456 ( .A(n163), .B(n23), .Z(SUM[9]) );
  COND1XL U457 ( .A(n164), .B(n166), .C(n165), .Z(n163) );
  CENX1 U458 ( .A(n174), .B(n25), .Z(SUM[7]) );
  COND1XL U459 ( .A(n175), .B(n177), .C(n176), .Z(n174) );
  CEOX1 U460 ( .A(n26), .B(n177), .Z(SUM[6]) );
  CEOX1 U461 ( .A(n27), .B(n182), .Z(SUM[5]) );
  CANR1XL U462 ( .A(n228), .B(n187), .C(n184), .Z(n182) );
  CNR2X1 U463 ( .A(A[30]), .B(B[30]), .Z(n34) );
  CNR2XL U464 ( .A(A[0]), .B(B[0]), .Z(n200) );
  CND2X1 U465 ( .A(A[29]), .B(B[29]), .Z(n40) );
  CND2X1 U466 ( .A(A[30]), .B(B[30]), .Z(n35) );
  COR2X1 U467 ( .A(A[29]), .B(B[29]), .Z(n338) );
  CENX1 U468 ( .A(n187), .B(n28), .Z(SUM[4]) );
  CENX1 U469 ( .A(n193), .B(n29), .Z(SUM[3]) );
  COND1XL U470 ( .A(n194), .B(n196), .C(n195), .Z(n193) );
  CEOX1 U471 ( .A(n30), .B(n196), .Z(SUM[2]) );
  CIVX2 U472 ( .A(n97), .Z(n95) );
  CIVX2 U473 ( .A(n94), .Z(n93) );
  CIVX2 U474 ( .A(n67), .Z(n69) );
  CIVX2 U475 ( .A(n60), .Z(n58) );
  CIVX2 U476 ( .A(n59), .Z(n57) );
  CIVX2 U477 ( .A(n48), .Z(n46) );
  CIVX2 U478 ( .A(n40), .Z(n38) );
  CIVX2 U479 ( .A(n198), .Z(n231) );
  CIVX2 U480 ( .A(n194), .Z(n230) );
  CIVX2 U481 ( .A(n191), .Z(n229) );
  CIVX2 U482 ( .A(n180), .Z(n227) );
  CIVX2 U483 ( .A(n175), .Z(n226) );
  CIVX2 U484 ( .A(n172), .Z(n225) );
  CIVX2 U485 ( .A(n164), .Z(n224) );
  CIVX2 U486 ( .A(n161), .Z(n223) );
  CIVX2 U487 ( .A(n149), .Z(n221) );
  CIVX2 U488 ( .A(n136), .Z(n219) );
  CIVX2 U489 ( .A(n124), .Z(n217) );
  CIVX2 U490 ( .A(n109), .Z(n215) );
  CIVX2 U491 ( .A(n104), .Z(n214) );
  CIVX2 U492 ( .A(n101), .Z(n213) );
  CIVX2 U493 ( .A(n91), .Z(n212) );
  CIVX2 U494 ( .A(n88), .Z(n211) );
  CIVX2 U495 ( .A(n83), .Z(n210) );
  CIVX2 U496 ( .A(n80), .Z(n209) );
  CIVX2 U497 ( .A(n66), .Z(n68) );
  CIVX2 U498 ( .A(n42), .Z(n204) );
  CIVX2 U499 ( .A(n34), .Z(n202) );
  CIVX2 U500 ( .A(n197), .Z(n196) );
  CIVX2 U501 ( .A(n188), .Z(n187) );
  CIVX2 U502 ( .A(n186), .Z(n184) );
  CIVX2 U503 ( .A(n167), .Z(n166) );
  CIVX2 U504 ( .A(n160), .Z(n158) );
  CIVX2 U505 ( .A(n159), .Z(n157) );
  CIVX2 U506 ( .A(n155), .Z(n153) );
  CIVX2 U507 ( .A(n154), .Z(n222) );
  CIVX2 U508 ( .A(n142), .Z(n140) );
  CIVX2 U509 ( .A(n141), .Z(n220) );
  CIVX2 U510 ( .A(n135), .Z(n133) );
  CIVX2 U511 ( .A(n134), .Z(n132) );
  CIVX2 U512 ( .A(n130), .Z(n128) );
  CIVX2 U513 ( .A(n129), .Z(n218) );
  CIVX2 U514 ( .A(n115), .Z(n113) );
  CIVX2 U515 ( .A(n114), .Z(n216) );
  CIVX2 U516 ( .A(n32), .Z(SUM[0]) );
endmodule


module calc_DW01_add_7 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n32, n33, n34, n35, n36, n38, n40, n41, n42, n43, n44, n46, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n187, n188, n190, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n326, n322, n323, n324, n325;

  CFA1X1 U3 ( .A(B[30]), .B(n33), .CI(A[30]), .CO(n32), .S(SUM[30]) );
  CAN2XL U252 ( .A(n323), .B(n187), .Z(SUM[0]) );
  CNIVX1 U253 ( .A(n326), .Z(SUM[1]) );
  CND2XL U254 ( .A(A[0]), .B(B[0]), .Z(n187) );
  COND1X2 U255 ( .A(n34), .B(n36), .C(n35), .Z(n33) );
  CANR1X2 U256 ( .A(n325), .B(n41), .C(n38), .Z(n36) );
  CANR1X2 U257 ( .A(n153), .B(n104), .C(n105), .Z(n103) );
  COND1X1 U258 ( .A(n154), .B(n174), .C(n155), .Z(n153) );
  COND1X1 U259 ( .A(n42), .B(n44), .C(n43), .Z(n41) );
  CND2XL U260 ( .A(A[6]), .B(B[6]), .Z(n162) );
  CNR2XL U261 ( .A(n161), .B(n158), .Z(n156) );
  CANR1XL U262 ( .A(n94), .B(n85), .C(n86), .Z(n84) );
  CANR1XL U263 ( .A(n52), .B(n61), .C(n53), .Z(n51) );
  COND1XL U264 ( .A(n187), .B(n184), .C(n185), .Z(n183) );
  CND2XL U265 ( .A(n216), .B(n185), .Z(n30) );
  CNR2X1 U266 ( .A(A[12]), .B(B[12]), .Z(n127) );
  CNR2XL U267 ( .A(n83), .B(n62), .Z(n60) );
  CIVX1 U268 ( .A(n80), .Z(n79) );
  COND1X1 U269 ( .A(n50), .B(n103), .C(n51), .Z(n49) );
  CND2XL U270 ( .A(n60), .B(n52), .Z(n50) );
  CND2XL U271 ( .A(n164), .B(n156), .Z(n154) );
  CNR2XL U272 ( .A(n127), .B(n122), .Z(n120) );
  CNR2XL U273 ( .A(n150), .B(n147), .Z(n145) );
  CNR2XL U274 ( .A(n90), .B(n87), .Z(n85) );
  CNR2XL U275 ( .A(n115), .B(n110), .Z(n108) );
  CNR2XL U276 ( .A(n140), .B(n135), .Z(n133) );
  CNR2XL U277 ( .A(n100), .B(n95), .Z(n93) );
  CEOXL U278 ( .A(n2), .B(n36), .Z(SUM[29]) );
  CND2XL U279 ( .A(n209), .B(n151), .Z(n23) );
  CND2XL U280 ( .A(n205), .B(n128), .Z(n19) );
  CND2XL U281 ( .A(n199), .B(n91), .Z(n13) );
  CEOXL U282 ( .A(n9), .B(n71), .Z(SUM[22]) );
  CEOXL U283 ( .A(n4), .B(n44), .Z(SUM[27]) );
  CND2XL U284 ( .A(n207), .B(n141), .Z(n21) );
  CND2XL U285 ( .A(n203), .B(n116), .Z(n17) );
  CND2XL U286 ( .A(n98), .B(n101), .Z(n15) );
  CND2XL U287 ( .A(n196), .B(n75), .Z(n10) );
  CEOXL U288 ( .A(n187), .B(n30), .Z(n326) );
  CND2XL U289 ( .A(n215), .B(n181), .Z(n29) );
  CND2XL U290 ( .A(n213), .B(n172), .Z(n27) );
  CNR2XL U291 ( .A(A[8]), .B(B[8]), .Z(n150) );
  CNR2XL U292 ( .A(A[16]), .B(B[16]), .Z(n100) );
  CENX1 U293 ( .A(n322), .B(n32), .Z(SUM[31]) );
  CENX1 U294 ( .A(B[31]), .B(A[31]), .Z(n322) );
  CND2XL U295 ( .A(A[20]), .B(B[20]), .Z(n78) );
  CND2XL U296 ( .A(A[22]), .B(B[22]), .Z(n70) );
  CND2XL U297 ( .A(A[24]), .B(B[24]), .Z(n58) );
  CND2XL U298 ( .A(A[1]), .B(B[1]), .Z(n185) );
  CND2XL U299 ( .A(A[3]), .B(B[3]), .Z(n178) );
  CND2XL U300 ( .A(A[9]), .B(B[9]), .Z(n148) );
  CND2XL U301 ( .A(A[13]), .B(B[13]), .Z(n123) );
  CND2XL U302 ( .A(A[7]), .B(B[7]), .Z(n159) );
  CND2XL U303 ( .A(A[5]), .B(B[5]), .Z(n167) );
  CND2XL U304 ( .A(A[11]), .B(B[11]), .Z(n136) );
  CND2XL U305 ( .A(A[15]), .B(B[15]), .Z(n111) );
  CND2XL U306 ( .A(A[19]), .B(B[19]), .Z(n88) );
  CND2XL U307 ( .A(A[17]), .B(B[17]), .Z(n96) );
  CND2XL U308 ( .A(A[23]), .B(B[23]), .Z(n67) );
  CND2XL U309 ( .A(A[25]), .B(B[25]), .Z(n55) );
  COR2XL U310 ( .A(A[0]), .B(B[0]), .Z(n323) );
  CANR1XL U311 ( .A(n164), .B(n173), .C(n165), .Z(n163) );
  CANR1XL U312 ( .A(n93), .B(n102), .C(n94), .Z(n92) );
  CANR1XL U313 ( .A(n72), .B(n79), .C(n73), .Z(n71) );
  CANR1XL U314 ( .A(n60), .B(n102), .C(n61), .Z(n59) );
  COND1XL U315 ( .A(n143), .B(n152), .C(n144), .Z(n142) );
  COND1XL U316 ( .A(n118), .B(n129), .C(n119), .Z(n117) );
  CNR2X1 U317 ( .A(n131), .B(n106), .Z(n104) );
  COND1XL U318 ( .A(n106), .B(n132), .C(n107), .Z(n105) );
  CND2X1 U319 ( .A(n120), .B(n108), .Z(n106) );
  CANR1XL U320 ( .A(n81), .B(n102), .C(n82), .Z(n80) );
  COND1XL U321 ( .A(n131), .B(n152), .C(n132), .Z(n130) );
  CND2X1 U322 ( .A(n93), .B(n85), .Z(n83) );
  CND2X1 U323 ( .A(n72), .B(n64), .Z(n62) );
  CND2X1 U324 ( .A(n145), .B(n133), .Z(n131) );
  CANR1XL U325 ( .A(n324), .B(n49), .C(n46), .Z(n44) );
  CNR2X1 U326 ( .A(n57), .B(n54), .Z(n52) );
  CENX1 U327 ( .A(n160), .B(n24), .Z(SUM[7]) );
  CND2X1 U328 ( .A(n210), .B(n159), .Z(n24) );
  COND1XL U329 ( .A(n161), .B(n163), .C(n162), .Z(n160) );
  CENX1 U330 ( .A(n68), .B(n8), .Z(SUM[23]) );
  CND2X1 U331 ( .A(n194), .B(n67), .Z(n8) );
  COND1XL U332 ( .A(n69), .B(n71), .C(n70), .Z(n68) );
  COND1XL U333 ( .A(n91), .B(n87), .C(n88), .Z(n86) );
  CANR1XL U334 ( .A(n183), .B(n175), .C(n176), .Z(n174) );
  CNR2X1 U335 ( .A(n180), .B(n177), .Z(n175) );
  COND1XL U336 ( .A(n181), .B(n177), .C(n178), .Z(n176) );
  CANR1XL U337 ( .A(n165), .B(n156), .C(n157), .Z(n155) );
  COND1XL U338 ( .A(n151), .B(n147), .C(n148), .Z(n146) );
  COND1XL U339 ( .A(n128), .B(n122), .C(n123), .Z(n121) );
  CANR1XL U340 ( .A(n146), .B(n133), .C(n134), .Z(n132) );
  COND1XL U341 ( .A(n141), .B(n135), .C(n136), .Z(n134) );
  COND1XL U342 ( .A(n172), .B(n166), .C(n167), .Z(n165) );
  COND1XL U343 ( .A(n101), .B(n95), .C(n96), .Z(n94) );
  COND1XL U344 ( .A(n78), .B(n74), .C(n75), .Z(n73) );
  COND1XL U345 ( .A(n62), .B(n84), .C(n63), .Z(n61) );
  CANR1XL U346 ( .A(n73), .B(n64), .C(n65), .Z(n63) );
  COND1XL U347 ( .A(n70), .B(n66), .C(n67), .Z(n65) );
  CANR1XL U348 ( .A(n121), .B(n108), .C(n109), .Z(n107) );
  COND1XL U349 ( .A(n116), .B(n110), .C(n111), .Z(n109) );
  CNR2X1 U350 ( .A(n69), .B(n66), .Z(n64) );
  CENX1 U351 ( .A(n149), .B(n22), .Z(SUM[9]) );
  CND2X1 U352 ( .A(n208), .B(n148), .Z(n22) );
  COND1XL U353 ( .A(n150), .B(n152), .C(n151), .Z(n149) );
  CENX1 U354 ( .A(n142), .B(n21), .Z(SUM[10]) );
  CENX1 U355 ( .A(n117), .B(n17), .Z(SUM[14]) );
  CENX1 U356 ( .A(n102), .B(n15), .Z(SUM[16]) );
  CENX1 U357 ( .A(n89), .B(n12), .Z(SUM[19]) );
  CND2X1 U358 ( .A(n198), .B(n88), .Z(n12) );
  COND1XL U359 ( .A(n90), .B(n92), .C(n91), .Z(n89) );
  CENX1 U360 ( .A(n79), .B(n11), .Z(SUM[20]) );
  CND2X1 U361 ( .A(n197), .B(n78), .Z(n11) );
  CENX1 U362 ( .A(n76), .B(n10), .Z(SUM[21]) );
  COND1XL U363 ( .A(n77), .B(n80), .C(n78), .Z(n76) );
  CENX1 U364 ( .A(n56), .B(n6), .Z(SUM[25]) );
  CND2X1 U365 ( .A(n192), .B(n55), .Z(n6) );
  COND1XL U366 ( .A(n57), .B(n59), .C(n58), .Z(n56) );
  CENX1 U367 ( .A(n49), .B(n5), .Z(SUM[26]) );
  CND2X1 U368 ( .A(n324), .B(n48), .Z(n5) );
  CENX1 U369 ( .A(n41), .B(n3), .Z(SUM[28]) );
  CND2X1 U370 ( .A(n325), .B(n40), .Z(n3) );
  COND1XL U371 ( .A(n162), .B(n158), .C(n159), .Z(n157) );
  COND1XL U372 ( .A(n58), .B(n54), .C(n55), .Z(n53) );
  CNR2X1 U373 ( .A(n171), .B(n166), .Z(n164) );
  CNR2X1 U374 ( .A(n77), .B(n74), .Z(n72) );
  CEOX1 U375 ( .A(n20), .B(n137), .Z(SUM[11]) );
  CND2X1 U376 ( .A(n206), .B(n136), .Z(n20) );
  CANR1XL U377 ( .A(n207), .B(n142), .C(n139), .Z(n137) );
  CEOX1 U378 ( .A(n19), .B(n129), .Z(SUM[12]) );
  CEOX1 U379 ( .A(n18), .B(n124), .Z(SUM[13]) );
  CND2X1 U380 ( .A(n204), .B(n123), .Z(n18) );
  CANR1XL U381 ( .A(n205), .B(n130), .C(n126), .Z(n124) );
  CEOX1 U382 ( .A(n16), .B(n112), .Z(SUM[15]) );
  CND2X1 U383 ( .A(n202), .B(n111), .Z(n16) );
  CANR1XL U384 ( .A(n203), .B(n117), .C(n114), .Z(n112) );
  CEOX1 U385 ( .A(n14), .B(n97), .Z(SUM[17]) );
  CND2X1 U386 ( .A(n200), .B(n96), .Z(n14) );
  CANR1XL U387 ( .A(n98), .B(n102), .C(n99), .Z(n97) );
  CEOX1 U388 ( .A(n13), .B(n92), .Z(SUM[18]) );
  CND2X1 U389 ( .A(n195), .B(n70), .Z(n9) );
  CEOX1 U390 ( .A(n7), .B(n59), .Z(SUM[24]) );
  CND2X1 U391 ( .A(n193), .B(n58), .Z(n7) );
  CND2X1 U392 ( .A(n190), .B(n43), .Z(n4) );
  CND2X1 U393 ( .A(n188), .B(n35), .Z(n2) );
  CEOX1 U394 ( .A(n26), .B(n168), .Z(SUM[5]) );
  CND2X1 U395 ( .A(n212), .B(n167), .Z(n26) );
  CANR1XL U396 ( .A(n213), .B(n173), .C(n170), .Z(n168) );
  CENX1 U397 ( .A(n179), .B(n28), .Z(SUM[3]) );
  CND2X1 U398 ( .A(n214), .B(n178), .Z(n28) );
  COND1XL U399 ( .A(n180), .B(n182), .C(n181), .Z(n179) );
  CENX1 U400 ( .A(n173), .B(n27), .Z(SUM[4]) );
  CEOX1 U401 ( .A(n29), .B(n182), .Z(SUM[2]) );
  CEOX1 U402 ( .A(n25), .B(n163), .Z(SUM[6]) );
  CND2X1 U403 ( .A(n211), .B(n162), .Z(n25) );
  CEOX1 U404 ( .A(n23), .B(n152), .Z(SUM[8]) );
  CNR2X1 U405 ( .A(A[5]), .B(B[5]), .Z(n166) );
  CNR2X1 U406 ( .A(A[17]), .B(B[17]), .Z(n95) );
  CNR2X1 U407 ( .A(A[19]), .B(B[19]), .Z(n87) );
  CNR2X1 U408 ( .A(A[21]), .B(B[21]), .Z(n74) );
  CNR2X1 U409 ( .A(A[23]), .B(B[23]), .Z(n66) );
  CNR2X1 U410 ( .A(A[9]), .B(B[9]), .Z(n147) );
  CNR2X1 U411 ( .A(A[3]), .B(B[3]), .Z(n177) );
  CNR2X1 U412 ( .A(A[11]), .B(B[11]), .Z(n135) );
  CNR2X1 U413 ( .A(A[15]), .B(B[15]), .Z(n110) );
  CNR2X1 U414 ( .A(A[13]), .B(B[13]), .Z(n122) );
  CNR2X1 U415 ( .A(A[7]), .B(B[7]), .Z(n158) );
  CNR2X1 U416 ( .A(A[25]), .B(B[25]), .Z(n54) );
  CNR2X1 U417 ( .A(A[2]), .B(B[2]), .Z(n180) );
  CNR2X1 U418 ( .A(A[6]), .B(B[6]), .Z(n161) );
  CNR2X1 U419 ( .A(A[18]), .B(B[18]), .Z(n90) );
  CNR2X1 U420 ( .A(A[20]), .B(B[20]), .Z(n77) );
  CNR2X1 U421 ( .A(A[22]), .B(B[22]), .Z(n69) );
  CNR2X1 U422 ( .A(A[24]), .B(B[24]), .Z(n57) );
  CNR2X1 U423 ( .A(A[14]), .B(B[14]), .Z(n115) );
  CNR2X1 U424 ( .A(A[10]), .B(B[10]), .Z(n140) );
  CNR2X1 U425 ( .A(A[4]), .B(B[4]), .Z(n171) );
  CNR2X1 U426 ( .A(A[27]), .B(B[27]), .Z(n42) );
  CNR2X1 U427 ( .A(A[1]), .B(B[1]), .Z(n184) );
  CND2X1 U428 ( .A(A[4]), .B(B[4]), .Z(n172) );
  CND2X1 U429 ( .A(A[10]), .B(B[10]), .Z(n141) );
  CND2X1 U430 ( .A(A[14]), .B(B[14]), .Z(n116) );
  CND2X1 U431 ( .A(A[12]), .B(B[12]), .Z(n128) );
  CND2X1 U432 ( .A(A[16]), .B(B[16]), .Z(n101) );
  CND2X1 U433 ( .A(A[2]), .B(B[2]), .Z(n181) );
  CND2X1 U434 ( .A(A[8]), .B(B[8]), .Z(n151) );
  CND2X1 U435 ( .A(A[18]), .B(B[18]), .Z(n91) );
  CND2X1 U436 ( .A(A[26]), .B(B[26]), .Z(n48) );
  CND2X1 U437 ( .A(A[28]), .B(B[28]), .Z(n40) );
  CND2X1 U438 ( .A(A[21]), .B(B[21]), .Z(n75) );
  CND2X1 U439 ( .A(A[27]), .B(B[27]), .Z(n43) );
  COR2X1 U440 ( .A(A[26]), .B(B[26]), .Z(n324) );
  COR2X1 U441 ( .A(A[28]), .B(B[28]), .Z(n325) );
  CNR2X1 U442 ( .A(A[29]), .B(B[29]), .Z(n34) );
  CND2X1 U443 ( .A(A[29]), .B(B[29]), .Z(n35) );
  CIVX2 U444 ( .A(n101), .Z(n99) );
  CIVX2 U445 ( .A(n84), .Z(n82) );
  CIVX2 U446 ( .A(n83), .Z(n81) );
  CIVX2 U447 ( .A(n48), .Z(n46) );
  CIVX2 U448 ( .A(n40), .Z(n38) );
  CIVX2 U449 ( .A(n184), .Z(n216) );
  CIVX2 U450 ( .A(n180), .Z(n215) );
  CIVX2 U451 ( .A(n177), .Z(n214) );
  CIVX2 U452 ( .A(n166), .Z(n212) );
  CIVX2 U453 ( .A(n161), .Z(n211) );
  CIVX2 U454 ( .A(n158), .Z(n210) );
  CIVX2 U455 ( .A(n150), .Z(n209) );
  CIVX2 U456 ( .A(n147), .Z(n208) );
  CIVX2 U457 ( .A(n135), .Z(n206) );
  CIVX2 U458 ( .A(n122), .Z(n204) );
  CIVX2 U459 ( .A(n110), .Z(n202) );
  CIVX2 U460 ( .A(n100), .Z(n98) );
  CIVX2 U461 ( .A(n95), .Z(n200) );
  CIVX2 U462 ( .A(n90), .Z(n199) );
  CIVX2 U463 ( .A(n87), .Z(n198) );
  CIVX2 U464 ( .A(n77), .Z(n197) );
  CIVX2 U465 ( .A(n74), .Z(n196) );
  CIVX2 U466 ( .A(n69), .Z(n195) );
  CIVX2 U467 ( .A(n66), .Z(n194) );
  CIVX2 U468 ( .A(n57), .Z(n193) );
  CIVX2 U469 ( .A(n54), .Z(n192) );
  CIVX2 U470 ( .A(n42), .Z(n190) );
  CIVX2 U471 ( .A(n34), .Z(n188) );
  CIVX2 U472 ( .A(n183), .Z(n182) );
  CIVX2 U473 ( .A(n174), .Z(n173) );
  CIVX2 U474 ( .A(n172), .Z(n170) );
  CIVX2 U475 ( .A(n171), .Z(n213) );
  CIVX2 U476 ( .A(n153), .Z(n152) );
  CIVX2 U477 ( .A(n146), .Z(n144) );
  CIVX2 U478 ( .A(n145), .Z(n143) );
  CIVX2 U479 ( .A(n141), .Z(n139) );
  CIVX2 U480 ( .A(n140), .Z(n207) );
  CIVX2 U481 ( .A(n130), .Z(n129) );
  CIVX2 U482 ( .A(n128), .Z(n126) );
  CIVX2 U483 ( .A(n127), .Z(n205) );
  CIVX2 U484 ( .A(n121), .Z(n119) );
  CIVX2 U485 ( .A(n120), .Z(n118) );
  CIVX2 U486 ( .A(n116), .Z(n114) );
  CIVX2 U487 ( .A(n115), .Z(n203) );
  CIVX2 U488 ( .A(n103), .Z(n102) );
endmodule


module calc_DW01_add_8 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n32, n33, n34, n35, n36, n38, n40, n41, n42, n43, n44, n46, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n187, n188, n190, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n326, n322, n323, n324, n325;

  CFA1X1 U3 ( .A(B[30]), .B(n33), .CI(A[30]), .CO(n32), .S(SUM[30]) );
  CAN2XL U252 ( .A(n322), .B(n187), .Z(SUM[0]) );
  CNIVX1 U253 ( .A(n326), .Z(SUM[1]) );
  CNR2XL U254 ( .A(A[1]), .B(B[1]), .Z(n184) );
  CANR1X1 U255 ( .A(n183), .B(n175), .C(n176), .Z(n174) );
  COND1X2 U256 ( .A(n34), .B(n36), .C(n35), .Z(n33) );
  CANR1X1 U257 ( .A(n325), .B(n41), .C(n38), .Z(n36) );
  CANR1X1 U258 ( .A(n153), .B(n104), .C(n105), .Z(n103) );
  COND1X1 U259 ( .A(n154), .B(n174), .C(n155), .Z(n153) );
  CND2XL U260 ( .A(A[6]), .B(B[6]), .Z(n162) );
  COND1XL U261 ( .A(n42), .B(n44), .C(n43), .Z(n41) );
  CNR2XL U262 ( .A(n161), .B(n158), .Z(n156) );
  CANR1XL U263 ( .A(n52), .B(n61), .C(n53), .Z(n51) );
  COND1XL U264 ( .A(n187), .B(n184), .C(n185), .Z(n183) );
  CND2XL U265 ( .A(n216), .B(n185), .Z(n30) );
  CNR2X1 U266 ( .A(A[12]), .B(B[12]), .Z(n127) );
  CNR2XL U267 ( .A(n83), .B(n62), .Z(n60) );
  CIVX1 U268 ( .A(n80), .Z(n79) );
  CIVXL U269 ( .A(n84), .Z(n82) );
  COND1X1 U270 ( .A(n50), .B(n103), .C(n51), .Z(n49) );
  CND2XL U271 ( .A(n60), .B(n52), .Z(n50) );
  CND2XL U272 ( .A(n164), .B(n156), .Z(n154) );
  CNR2XL U273 ( .A(n127), .B(n122), .Z(n120) );
  CNR2XL U274 ( .A(n150), .B(n147), .Z(n145) );
  CNR2XL U275 ( .A(n90), .B(n87), .Z(n85) );
  CNR2XL U276 ( .A(n115), .B(n110), .Z(n108) );
  CNR2XL U277 ( .A(n140), .B(n135), .Z(n133) );
  CNR2XL U278 ( .A(n100), .B(n95), .Z(n93) );
  CEOXL U279 ( .A(n2), .B(n36), .Z(SUM[29]) );
  CND2XL U280 ( .A(n209), .B(n151), .Z(n23) );
  CND2XL U281 ( .A(n205), .B(n128), .Z(n19) );
  CND2XL U282 ( .A(n199), .B(n91), .Z(n13) );
  CND2XL U283 ( .A(n195), .B(n70), .Z(n9) );
  CEOXL U284 ( .A(n9), .B(n71), .Z(SUM[22]) );
  CEOXL U285 ( .A(n4), .B(n44), .Z(SUM[27]) );
  CND2XL U286 ( .A(n194), .B(n67), .Z(n8) );
  CND2XL U287 ( .A(n207), .B(n141), .Z(n21) );
  CND2XL U288 ( .A(n203), .B(n116), .Z(n17) );
  CND2XL U289 ( .A(n98), .B(n101), .Z(n15) );
  CND2XL U290 ( .A(n197), .B(n78), .Z(n11) );
  CND2XL U291 ( .A(n196), .B(n75), .Z(n10) );
  CEOXL U292 ( .A(n187), .B(n30), .Z(n326) );
  CND2XL U293 ( .A(n215), .B(n181), .Z(n29) );
  CND2XL U294 ( .A(n213), .B(n172), .Z(n27) );
  CNR2XL U295 ( .A(A[8]), .B(B[8]), .Z(n150) );
  CNR2XL U296 ( .A(A[16]), .B(B[16]), .Z(n100) );
  CND2XL U297 ( .A(A[1]), .B(B[1]), .Z(n185) );
  CND2XL U298 ( .A(A[3]), .B(B[3]), .Z(n178) );
  CND2XL U299 ( .A(A[9]), .B(B[9]), .Z(n148) );
  CND2XL U300 ( .A(A[13]), .B(B[13]), .Z(n123) );
  CND2XL U301 ( .A(A[7]), .B(B[7]), .Z(n159) );
  CND2XL U302 ( .A(A[5]), .B(B[5]), .Z(n167) );
  CND2XL U303 ( .A(A[11]), .B(B[11]), .Z(n136) );
  CND2XL U304 ( .A(A[15]), .B(B[15]), .Z(n111) );
  CND2XL U305 ( .A(A[19]), .B(B[19]), .Z(n88) );
  CND2XL U306 ( .A(A[17]), .B(B[17]), .Z(n96) );
  COR2XL U307 ( .A(A[0]), .B(B[0]), .Z(n322) );
  CANR1XL U308 ( .A(n164), .B(n173), .C(n165), .Z(n163) );
  CANR1XL U309 ( .A(n93), .B(n102), .C(n94), .Z(n92) );
  CANR1XL U310 ( .A(n72), .B(n79), .C(n73), .Z(n71) );
  CANR1XL U311 ( .A(n60), .B(n102), .C(n61), .Z(n59) );
  COND1XL U312 ( .A(n143), .B(n152), .C(n144), .Z(n142) );
  COND1XL U313 ( .A(n118), .B(n129), .C(n119), .Z(n117) );
  CNR2X1 U314 ( .A(n131), .B(n106), .Z(n104) );
  COND1XL U315 ( .A(n106), .B(n132), .C(n107), .Z(n105) );
  CND2X1 U316 ( .A(n120), .B(n108), .Z(n106) );
  CANR1XL U317 ( .A(n81), .B(n102), .C(n82), .Z(n80) );
  COND1XL U318 ( .A(n131), .B(n152), .C(n132), .Z(n130) );
  CND2X1 U319 ( .A(n93), .B(n85), .Z(n83) );
  CND2X1 U320 ( .A(n72), .B(n64), .Z(n62) );
  CND2X1 U321 ( .A(n145), .B(n133), .Z(n131) );
  CANR1XL U322 ( .A(n324), .B(n49), .C(n46), .Z(n44) );
  CNR2X1 U323 ( .A(n57), .B(n54), .Z(n52) );
  CENX1 U324 ( .A(n160), .B(n24), .Z(SUM[7]) );
  CND2X1 U325 ( .A(n210), .B(n159), .Z(n24) );
  COND1XL U326 ( .A(n161), .B(n163), .C(n162), .Z(n160) );
  CENX1 U327 ( .A(n68), .B(n8), .Z(SUM[23]) );
  COND1XL U328 ( .A(n69), .B(n71), .C(n70), .Z(n68) );
  CANR1XL U329 ( .A(n94), .B(n85), .C(n86), .Z(n84) );
  COND1XL U330 ( .A(n91), .B(n87), .C(n88), .Z(n86) );
  CNR2X1 U331 ( .A(n180), .B(n177), .Z(n175) );
  COND1XL U332 ( .A(n181), .B(n177), .C(n178), .Z(n176) );
  CANR1XL U333 ( .A(n165), .B(n156), .C(n157), .Z(n155) );
  COND1XL U334 ( .A(n151), .B(n147), .C(n148), .Z(n146) );
  COND1XL U335 ( .A(n128), .B(n122), .C(n123), .Z(n121) );
  CANR1XL U336 ( .A(n146), .B(n133), .C(n134), .Z(n132) );
  COND1XL U337 ( .A(n141), .B(n135), .C(n136), .Z(n134) );
  COND1XL U338 ( .A(n172), .B(n166), .C(n167), .Z(n165) );
  COND1XL U339 ( .A(n101), .B(n95), .C(n96), .Z(n94) );
  COND1XL U340 ( .A(n78), .B(n74), .C(n75), .Z(n73) );
  COND1XL U341 ( .A(n62), .B(n84), .C(n63), .Z(n61) );
  CANR1XL U342 ( .A(n73), .B(n64), .C(n65), .Z(n63) );
  COND1XL U343 ( .A(n70), .B(n66), .C(n67), .Z(n65) );
  CANR1XL U344 ( .A(n121), .B(n108), .C(n109), .Z(n107) );
  COND1XL U345 ( .A(n116), .B(n110), .C(n111), .Z(n109) );
  CNR2X1 U346 ( .A(n69), .B(n66), .Z(n64) );
  CENX1 U347 ( .A(n149), .B(n22), .Z(SUM[9]) );
  CND2X1 U348 ( .A(n208), .B(n148), .Z(n22) );
  COND1XL U349 ( .A(n150), .B(n152), .C(n151), .Z(n149) );
  CENX1 U350 ( .A(n142), .B(n21), .Z(SUM[10]) );
  CENX1 U351 ( .A(n117), .B(n17), .Z(SUM[14]) );
  CENX1 U352 ( .A(n102), .B(n15), .Z(SUM[16]) );
  CENX1 U353 ( .A(n89), .B(n12), .Z(SUM[19]) );
  CND2X1 U354 ( .A(n198), .B(n88), .Z(n12) );
  COND1XL U355 ( .A(n90), .B(n92), .C(n91), .Z(n89) );
  CENX1 U356 ( .A(n79), .B(n11), .Z(SUM[20]) );
  CENX1 U357 ( .A(n76), .B(n10), .Z(SUM[21]) );
  COND1XL U358 ( .A(n77), .B(n80), .C(n78), .Z(n76) );
  CENX1 U359 ( .A(n56), .B(n6), .Z(SUM[25]) );
  CND2X1 U360 ( .A(n192), .B(n55), .Z(n6) );
  COND1XL U361 ( .A(n57), .B(n59), .C(n58), .Z(n56) );
  CENX1 U362 ( .A(n49), .B(n5), .Z(SUM[26]) );
  CND2X1 U363 ( .A(n324), .B(n48), .Z(n5) );
  CENX1 U364 ( .A(n41), .B(n3), .Z(SUM[28]) );
  CND2X1 U365 ( .A(n325), .B(n40), .Z(n3) );
  COND1XL U366 ( .A(n162), .B(n158), .C(n159), .Z(n157) );
  COND1XL U367 ( .A(n58), .B(n54), .C(n55), .Z(n53) );
  CNR2X1 U368 ( .A(n171), .B(n166), .Z(n164) );
  CNR2X1 U369 ( .A(n77), .B(n74), .Z(n72) );
  CEOX1 U370 ( .A(n20), .B(n137), .Z(SUM[11]) );
  CND2X1 U371 ( .A(n206), .B(n136), .Z(n20) );
  CANR1XL U372 ( .A(n207), .B(n142), .C(n139), .Z(n137) );
  CEOX1 U373 ( .A(n19), .B(n129), .Z(SUM[12]) );
  CEOX1 U374 ( .A(n18), .B(n124), .Z(SUM[13]) );
  CND2X1 U375 ( .A(n204), .B(n123), .Z(n18) );
  CANR1XL U376 ( .A(n205), .B(n130), .C(n126), .Z(n124) );
  CEOX1 U377 ( .A(n16), .B(n112), .Z(SUM[15]) );
  CND2X1 U378 ( .A(n202), .B(n111), .Z(n16) );
  CANR1XL U379 ( .A(n203), .B(n117), .C(n114), .Z(n112) );
  CEOX1 U380 ( .A(n14), .B(n97), .Z(SUM[17]) );
  CND2X1 U381 ( .A(n200), .B(n96), .Z(n14) );
  CANR1XL U382 ( .A(n98), .B(n102), .C(n99), .Z(n97) );
  CEOX1 U383 ( .A(n13), .B(n92), .Z(SUM[18]) );
  CEOX1 U384 ( .A(n7), .B(n59), .Z(SUM[24]) );
  CND2X1 U385 ( .A(n193), .B(n58), .Z(n7) );
  CND2X1 U386 ( .A(n190), .B(n43), .Z(n4) );
  CND2X1 U387 ( .A(n188), .B(n35), .Z(n2) );
  CEOX1 U388 ( .A(n26), .B(n168), .Z(SUM[5]) );
  CND2X1 U389 ( .A(n212), .B(n167), .Z(n26) );
  CANR1XL U390 ( .A(n213), .B(n173), .C(n170), .Z(n168) );
  CENX1 U391 ( .A(n179), .B(n28), .Z(SUM[3]) );
  CND2X1 U392 ( .A(n214), .B(n178), .Z(n28) );
  COND1XL U393 ( .A(n180), .B(n182), .C(n181), .Z(n179) );
  CENX1 U394 ( .A(n173), .B(n27), .Z(SUM[4]) );
  CEOX1 U395 ( .A(n29), .B(n182), .Z(SUM[2]) );
  CEOX1 U396 ( .A(n25), .B(n163), .Z(SUM[6]) );
  CND2X1 U397 ( .A(n211), .B(n162), .Z(n25) );
  CEOX1 U398 ( .A(n23), .B(n152), .Z(SUM[8]) );
  CNR2X1 U399 ( .A(A[5]), .B(B[5]), .Z(n166) );
  CNR2X1 U400 ( .A(A[17]), .B(B[17]), .Z(n95) );
  CNR2X1 U401 ( .A(A[19]), .B(B[19]), .Z(n87) );
  CNR2X1 U402 ( .A(A[21]), .B(B[21]), .Z(n74) );
  CNR2X1 U403 ( .A(A[23]), .B(B[23]), .Z(n66) );
  CNR2X1 U404 ( .A(A[9]), .B(B[9]), .Z(n147) );
  CNR2X1 U405 ( .A(A[3]), .B(B[3]), .Z(n177) );
  CNR2X1 U406 ( .A(A[11]), .B(B[11]), .Z(n135) );
  CNR2X1 U407 ( .A(A[15]), .B(B[15]), .Z(n110) );
  CNR2X1 U408 ( .A(A[13]), .B(B[13]), .Z(n122) );
  CNR2X1 U409 ( .A(A[7]), .B(B[7]), .Z(n158) );
  CNR2X1 U410 ( .A(A[25]), .B(B[25]), .Z(n54) );
  CNR2X1 U411 ( .A(A[2]), .B(B[2]), .Z(n180) );
  CNR2X1 U412 ( .A(A[6]), .B(B[6]), .Z(n161) );
  CNR2X1 U413 ( .A(A[18]), .B(B[18]), .Z(n90) );
  CNR2X1 U414 ( .A(A[20]), .B(B[20]), .Z(n77) );
  CNR2X1 U415 ( .A(A[22]), .B(B[22]), .Z(n69) );
  CNR2X1 U416 ( .A(A[24]), .B(B[24]), .Z(n57) );
  CNR2X1 U417 ( .A(A[14]), .B(B[14]), .Z(n115) );
  CNR2X1 U418 ( .A(A[10]), .B(B[10]), .Z(n140) );
  CNR2X1 U419 ( .A(A[4]), .B(B[4]), .Z(n171) );
  CND2X1 U420 ( .A(A[0]), .B(B[0]), .Z(n187) );
  CNR2X1 U421 ( .A(A[27]), .B(B[27]), .Z(n42) );
  CENX1 U422 ( .A(n323), .B(n32), .Z(SUM[31]) );
  CENX1 U423 ( .A(B[31]), .B(A[31]), .Z(n323) );
  CND2X1 U424 ( .A(A[4]), .B(B[4]), .Z(n172) );
  CND2X1 U425 ( .A(A[10]), .B(B[10]), .Z(n141) );
  CND2X1 U426 ( .A(A[14]), .B(B[14]), .Z(n116) );
  CND2X1 U427 ( .A(A[12]), .B(B[12]), .Z(n128) );
  CND2X1 U428 ( .A(A[16]), .B(B[16]), .Z(n101) );
  CND2X1 U429 ( .A(A[2]), .B(B[2]), .Z(n181) );
  CND2X1 U430 ( .A(A[8]), .B(B[8]), .Z(n151) );
  CND2X1 U431 ( .A(A[18]), .B(B[18]), .Z(n91) );
  CND2X1 U432 ( .A(A[20]), .B(B[20]), .Z(n78) );
  CND2X1 U433 ( .A(A[22]), .B(B[22]), .Z(n70) );
  CND2X1 U434 ( .A(A[24]), .B(B[24]), .Z(n58) );
  CND2X1 U435 ( .A(A[26]), .B(B[26]), .Z(n48) );
  CND2X1 U436 ( .A(A[28]), .B(B[28]), .Z(n40) );
  CND2X1 U437 ( .A(A[21]), .B(B[21]), .Z(n75) );
  CND2X1 U438 ( .A(A[23]), .B(B[23]), .Z(n67) );
  CND2X1 U439 ( .A(A[27]), .B(B[27]), .Z(n43) );
  CND2X1 U440 ( .A(A[25]), .B(B[25]), .Z(n55) );
  COR2X1 U441 ( .A(A[26]), .B(B[26]), .Z(n324) );
  COR2X1 U442 ( .A(A[28]), .B(B[28]), .Z(n325) );
  CNR2X1 U443 ( .A(A[29]), .B(B[29]), .Z(n34) );
  CND2X1 U444 ( .A(A[29]), .B(B[29]), .Z(n35) );
  CIVX2 U445 ( .A(n101), .Z(n99) );
  CIVX2 U446 ( .A(n83), .Z(n81) );
  CIVX2 U447 ( .A(n48), .Z(n46) );
  CIVX2 U448 ( .A(n40), .Z(n38) );
  CIVX2 U449 ( .A(n184), .Z(n216) );
  CIVX2 U450 ( .A(n180), .Z(n215) );
  CIVX2 U451 ( .A(n177), .Z(n214) );
  CIVX2 U452 ( .A(n166), .Z(n212) );
  CIVX2 U453 ( .A(n161), .Z(n211) );
  CIVX2 U454 ( .A(n158), .Z(n210) );
  CIVX2 U455 ( .A(n150), .Z(n209) );
  CIVX2 U456 ( .A(n147), .Z(n208) );
  CIVX2 U457 ( .A(n135), .Z(n206) );
  CIVX2 U458 ( .A(n122), .Z(n204) );
  CIVX2 U459 ( .A(n110), .Z(n202) );
  CIVX2 U460 ( .A(n100), .Z(n98) );
  CIVX2 U461 ( .A(n95), .Z(n200) );
  CIVX2 U462 ( .A(n90), .Z(n199) );
  CIVX2 U463 ( .A(n87), .Z(n198) );
  CIVX2 U464 ( .A(n77), .Z(n197) );
  CIVX2 U465 ( .A(n74), .Z(n196) );
  CIVX2 U466 ( .A(n69), .Z(n195) );
  CIVX2 U467 ( .A(n66), .Z(n194) );
  CIVX2 U468 ( .A(n57), .Z(n193) );
  CIVX2 U469 ( .A(n54), .Z(n192) );
  CIVX2 U470 ( .A(n42), .Z(n190) );
  CIVX2 U471 ( .A(n34), .Z(n188) );
  CIVX2 U472 ( .A(n183), .Z(n182) );
  CIVX2 U473 ( .A(n174), .Z(n173) );
  CIVX2 U474 ( .A(n172), .Z(n170) );
  CIVX2 U475 ( .A(n171), .Z(n213) );
  CIVX2 U476 ( .A(n153), .Z(n152) );
  CIVX2 U477 ( .A(n146), .Z(n144) );
  CIVX2 U478 ( .A(n145), .Z(n143) );
  CIVX2 U479 ( .A(n141), .Z(n139) );
  CIVX2 U480 ( .A(n140), .Z(n207) );
  CIVX2 U481 ( .A(n130), .Z(n129) );
  CIVX2 U482 ( .A(n128), .Z(n126) );
  CIVX2 U483 ( .A(n127), .Z(n205) );
  CIVX2 U484 ( .A(n121), .Z(n119) );
  CIVX2 U485 ( .A(n120), .Z(n118) );
  CIVX2 U486 ( .A(n116), .Z(n114) );
  CIVX2 U487 ( .A(n115), .Z(n203) );
  CIVX2 U488 ( .A(n103), .Z(n102) );
endmodule


module calc_DW01_add_9 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n32, n33, n34, n35, n36, n38, n40, n41, n42, n43, n44, n46, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n187,
         n188, n190, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n326, n322, n323, n324, n325;

  CFA1X1 U3 ( .A(B[30]), .B(n33), .CI(A[30]), .CO(n32), .S(SUM[30]) );
  CIVX2 U252 ( .A(n216), .Z(n30) );
  CNR2X2 U253 ( .A(n187), .B(n184), .Z(n183) );
  CIVX2 U254 ( .A(A[1]), .Z(n184) );
  CAN2XL U255 ( .A(n322), .B(n187), .Z(SUM[0]) );
  CNIVX1 U256 ( .A(n326), .Z(SUM[1]) );
  CND2XL U257 ( .A(A[0]), .B(B[0]), .Z(n187) );
  COND1X2 U258 ( .A(n34), .B(n36), .C(n35), .Z(n33) );
  CANR1X2 U259 ( .A(n325), .B(n41), .C(n38), .Z(n36) );
  CANR1X1 U260 ( .A(n153), .B(n104), .C(n105), .Z(n103) );
  COND1X1 U261 ( .A(n154), .B(n174), .C(n155), .Z(n153) );
  COND1X1 U262 ( .A(n42), .B(n44), .C(n43), .Z(n41) );
  CND2XL U263 ( .A(A[6]), .B(B[6]), .Z(n162) );
  CNR2XL U264 ( .A(n161), .B(n158), .Z(n156) );
  CANR1XL U265 ( .A(n52), .B(n61), .C(n53), .Z(n51) );
  CNR2X1 U266 ( .A(A[12]), .B(B[12]), .Z(n127) );
  CNR2XL U267 ( .A(n83), .B(n62), .Z(n60) );
  CIVX1 U268 ( .A(n80), .Z(n79) );
  CIVXL U269 ( .A(n84), .Z(n82) );
  COND1X1 U270 ( .A(n50), .B(n103), .C(n51), .Z(n49) );
  CND2XL U271 ( .A(n60), .B(n52), .Z(n50) );
  CND2XL U272 ( .A(n164), .B(n156), .Z(n154) );
  CNR2XL U273 ( .A(n127), .B(n122), .Z(n120) );
  CNR2XL U274 ( .A(n150), .B(n147), .Z(n145) );
  CNR2XL U275 ( .A(n90), .B(n87), .Z(n85) );
  CNR2XL U276 ( .A(n115), .B(n110), .Z(n108) );
  CNR2XL U277 ( .A(n140), .B(n135), .Z(n133) );
  CNR2XL U278 ( .A(n100), .B(n95), .Z(n93) );
  CEOXL U279 ( .A(n2), .B(n36), .Z(SUM[29]) );
  CND2XL U280 ( .A(n209), .B(n151), .Z(n23) );
  CND2XL U281 ( .A(n205), .B(n128), .Z(n19) );
  CND2XL U282 ( .A(n199), .B(n91), .Z(n13) );
  CND2XL U283 ( .A(n195), .B(n70), .Z(n9) );
  CEOXL U284 ( .A(n9), .B(n71), .Z(SUM[22]) );
  CEOXL U285 ( .A(n4), .B(n44), .Z(SUM[27]) );
  CND2XL U286 ( .A(n194), .B(n67), .Z(n8) );
  CND2XL U287 ( .A(n207), .B(n141), .Z(n21) );
  CND2XL U288 ( .A(n203), .B(n116), .Z(n17) );
  CND2XL U289 ( .A(n98), .B(n101), .Z(n15) );
  CND2XL U290 ( .A(n197), .B(n78), .Z(n11) );
  CND2XL U291 ( .A(n196), .B(n75), .Z(n10) );
  CND2XL U292 ( .A(n215), .B(n181), .Z(n29) );
  CND2XL U293 ( .A(n213), .B(n172), .Z(n27) );
  CNR2XL U294 ( .A(A[8]), .B(B[8]), .Z(n150) );
  CNR2XL U295 ( .A(A[16]), .B(B[16]), .Z(n100) );
  CND2XL U296 ( .A(A[3]), .B(B[3]), .Z(n178) );
  CND2XL U297 ( .A(A[9]), .B(B[9]), .Z(n148) );
  CND2XL U298 ( .A(A[13]), .B(B[13]), .Z(n123) );
  CND2XL U299 ( .A(A[7]), .B(B[7]), .Z(n159) );
  CND2XL U300 ( .A(A[5]), .B(B[5]), .Z(n167) );
  CND2XL U301 ( .A(A[11]), .B(B[11]), .Z(n136) );
  CND2XL U302 ( .A(A[15]), .B(B[15]), .Z(n111) );
  CND2XL U303 ( .A(A[19]), .B(B[19]), .Z(n88) );
  CND2XL U304 ( .A(A[17]), .B(B[17]), .Z(n96) );
  COR2XL U305 ( .A(A[0]), .B(B[0]), .Z(n322) );
  CANR1XL U306 ( .A(n164), .B(n173), .C(n165), .Z(n163) );
  CANR1XL U307 ( .A(n93), .B(n102), .C(n94), .Z(n92) );
  CANR1XL U308 ( .A(n72), .B(n79), .C(n73), .Z(n71) );
  CANR1XL U309 ( .A(n60), .B(n102), .C(n61), .Z(n59) );
  COND1XL U310 ( .A(n143), .B(n152), .C(n144), .Z(n142) );
  COND1XL U311 ( .A(n118), .B(n129), .C(n119), .Z(n117) );
  CNR2X1 U312 ( .A(n131), .B(n106), .Z(n104) );
  COND1XL U313 ( .A(n106), .B(n132), .C(n107), .Z(n105) );
  CND2X1 U314 ( .A(n120), .B(n108), .Z(n106) );
  CANR1XL U315 ( .A(n81), .B(n102), .C(n82), .Z(n80) );
  COND1XL U316 ( .A(n131), .B(n152), .C(n132), .Z(n130) );
  CND2X1 U317 ( .A(n93), .B(n85), .Z(n83) );
  CND2X1 U318 ( .A(n72), .B(n64), .Z(n62) );
  CND2X1 U319 ( .A(n145), .B(n133), .Z(n131) );
  CANR1XL U320 ( .A(n324), .B(n49), .C(n46), .Z(n44) );
  CNR2X1 U321 ( .A(n57), .B(n54), .Z(n52) );
  CENX1 U322 ( .A(n160), .B(n24), .Z(SUM[7]) );
  CND2X1 U323 ( .A(n210), .B(n159), .Z(n24) );
  COND1XL U324 ( .A(n161), .B(n163), .C(n162), .Z(n160) );
  CENX1 U325 ( .A(n68), .B(n8), .Z(SUM[23]) );
  COND1XL U326 ( .A(n69), .B(n71), .C(n70), .Z(n68) );
  CANR1XL U327 ( .A(n94), .B(n85), .C(n86), .Z(n84) );
  COND1XL U328 ( .A(n91), .B(n87), .C(n88), .Z(n86) );
  CANR1XL U329 ( .A(n183), .B(n175), .C(n176), .Z(n174) );
  CNR2X1 U330 ( .A(n180), .B(n177), .Z(n175) );
  COND1XL U331 ( .A(n181), .B(n177), .C(n178), .Z(n176) );
  CANR1XL U332 ( .A(n165), .B(n156), .C(n157), .Z(n155) );
  COND1XL U333 ( .A(n151), .B(n147), .C(n148), .Z(n146) );
  COND1XL U334 ( .A(n128), .B(n122), .C(n123), .Z(n121) );
  CANR1XL U335 ( .A(n146), .B(n133), .C(n134), .Z(n132) );
  COND1XL U336 ( .A(n141), .B(n135), .C(n136), .Z(n134) );
  COND1XL U337 ( .A(n172), .B(n166), .C(n167), .Z(n165) );
  COND1XL U338 ( .A(n101), .B(n95), .C(n96), .Z(n94) );
  COND1XL U339 ( .A(n78), .B(n74), .C(n75), .Z(n73) );
  COND1XL U340 ( .A(n62), .B(n84), .C(n63), .Z(n61) );
  CANR1XL U341 ( .A(n73), .B(n64), .C(n65), .Z(n63) );
  COND1XL U342 ( .A(n70), .B(n66), .C(n67), .Z(n65) );
  CANR1XL U343 ( .A(n121), .B(n108), .C(n109), .Z(n107) );
  COND1XL U344 ( .A(n116), .B(n110), .C(n111), .Z(n109) );
  CNR2X1 U345 ( .A(n69), .B(n66), .Z(n64) );
  CENX1 U346 ( .A(n149), .B(n22), .Z(SUM[9]) );
  CND2X1 U347 ( .A(n208), .B(n148), .Z(n22) );
  COND1XL U348 ( .A(n150), .B(n152), .C(n151), .Z(n149) );
  CENX1 U349 ( .A(n142), .B(n21), .Z(SUM[10]) );
  CENX1 U350 ( .A(n117), .B(n17), .Z(SUM[14]) );
  CENX1 U351 ( .A(n102), .B(n15), .Z(SUM[16]) );
  CENX1 U352 ( .A(n89), .B(n12), .Z(SUM[19]) );
  CND2X1 U353 ( .A(n198), .B(n88), .Z(n12) );
  COND1XL U354 ( .A(n90), .B(n92), .C(n91), .Z(n89) );
  CENX1 U355 ( .A(n79), .B(n11), .Z(SUM[20]) );
  CENX1 U356 ( .A(n76), .B(n10), .Z(SUM[21]) );
  COND1XL U357 ( .A(n77), .B(n80), .C(n78), .Z(n76) );
  CENX1 U358 ( .A(n56), .B(n6), .Z(SUM[25]) );
  CND2X1 U359 ( .A(n192), .B(n55), .Z(n6) );
  COND1XL U360 ( .A(n57), .B(n59), .C(n58), .Z(n56) );
  CENX1 U361 ( .A(n49), .B(n5), .Z(SUM[26]) );
  CND2X1 U362 ( .A(n324), .B(n48), .Z(n5) );
  CENX1 U363 ( .A(n41), .B(n3), .Z(SUM[28]) );
  CND2X1 U364 ( .A(n325), .B(n40), .Z(n3) );
  COND1XL U365 ( .A(n162), .B(n158), .C(n159), .Z(n157) );
  COND1XL U366 ( .A(n58), .B(n54), .C(n55), .Z(n53) );
  CNR2X1 U367 ( .A(n171), .B(n166), .Z(n164) );
  CNR2X1 U368 ( .A(n77), .B(n74), .Z(n72) );
  CEOX1 U369 ( .A(n20), .B(n137), .Z(SUM[11]) );
  CND2X1 U370 ( .A(n206), .B(n136), .Z(n20) );
  CANR1XL U371 ( .A(n207), .B(n142), .C(n139), .Z(n137) );
  CEOX1 U372 ( .A(n19), .B(n129), .Z(SUM[12]) );
  CEOX1 U373 ( .A(n18), .B(n124), .Z(SUM[13]) );
  CND2X1 U374 ( .A(n204), .B(n123), .Z(n18) );
  CANR1XL U375 ( .A(n205), .B(n130), .C(n126), .Z(n124) );
  CEOX1 U376 ( .A(n16), .B(n112), .Z(SUM[15]) );
  CND2X1 U377 ( .A(n202), .B(n111), .Z(n16) );
  CANR1XL U378 ( .A(n203), .B(n117), .C(n114), .Z(n112) );
  CEOX1 U379 ( .A(n14), .B(n97), .Z(SUM[17]) );
  CND2X1 U380 ( .A(n200), .B(n96), .Z(n14) );
  CANR1XL U381 ( .A(n98), .B(n102), .C(n99), .Z(n97) );
  CEOX1 U382 ( .A(n13), .B(n92), .Z(SUM[18]) );
  CEOX1 U383 ( .A(n7), .B(n59), .Z(SUM[24]) );
  CND2X1 U384 ( .A(n193), .B(n58), .Z(n7) );
  CND2X1 U385 ( .A(n190), .B(n43), .Z(n4) );
  CND2X1 U386 ( .A(n188), .B(n35), .Z(n2) );
  CEOX1 U387 ( .A(n26), .B(n168), .Z(SUM[5]) );
  CND2X1 U388 ( .A(n212), .B(n167), .Z(n26) );
  CANR1XL U389 ( .A(n213), .B(n173), .C(n170), .Z(n168) );
  CENX1 U390 ( .A(n179), .B(n28), .Z(SUM[3]) );
  CND2X1 U391 ( .A(n214), .B(n178), .Z(n28) );
  COND1XL U392 ( .A(n180), .B(n182), .C(n181), .Z(n179) );
  CENX1 U393 ( .A(n173), .B(n27), .Z(SUM[4]) );
  CEOX1 U394 ( .A(n29), .B(n182), .Z(SUM[2]) );
  CEOX1 U395 ( .A(n25), .B(n163), .Z(SUM[6]) );
  CND2X1 U396 ( .A(n211), .B(n162), .Z(n25) );
  CEOX1 U397 ( .A(n23), .B(n152), .Z(SUM[8]) );
  CNR2X1 U398 ( .A(A[5]), .B(B[5]), .Z(n166) );
  CNR2X1 U399 ( .A(A[17]), .B(B[17]), .Z(n95) );
  CNR2X1 U400 ( .A(A[19]), .B(B[19]), .Z(n87) );
  CNR2X1 U401 ( .A(A[21]), .B(B[21]), .Z(n74) );
  CNR2X1 U402 ( .A(A[23]), .B(B[23]), .Z(n66) );
  CNR2X1 U403 ( .A(A[9]), .B(B[9]), .Z(n147) );
  CNR2X1 U404 ( .A(A[3]), .B(B[3]), .Z(n177) );
  CNR2X1 U405 ( .A(A[11]), .B(B[11]), .Z(n135) );
  CNR2X1 U406 ( .A(A[15]), .B(B[15]), .Z(n110) );
  CNR2X1 U407 ( .A(A[13]), .B(B[13]), .Z(n122) );
  CNR2X1 U408 ( .A(A[7]), .B(B[7]), .Z(n158) );
  CNR2X1 U409 ( .A(A[25]), .B(B[25]), .Z(n54) );
  CNR2X1 U410 ( .A(A[2]), .B(B[2]), .Z(n180) );
  CNR2X1 U411 ( .A(A[6]), .B(B[6]), .Z(n161) );
  CNR2X1 U412 ( .A(A[18]), .B(B[18]), .Z(n90) );
  CNR2X1 U413 ( .A(A[20]), .B(B[20]), .Z(n77) );
  CNR2X1 U414 ( .A(A[22]), .B(B[22]), .Z(n69) );
  CNR2X1 U415 ( .A(A[24]), .B(B[24]), .Z(n57) );
  CNR2X1 U416 ( .A(A[14]), .B(B[14]), .Z(n115) );
  CNR2X1 U417 ( .A(A[10]), .B(B[10]), .Z(n140) );
  CNR2X1 U418 ( .A(A[4]), .B(B[4]), .Z(n171) );
  CNR2X1 U419 ( .A(A[27]), .B(B[27]), .Z(n42) );
  CENX1 U420 ( .A(n323), .B(n32), .Z(SUM[31]) );
  CENX1 U421 ( .A(B[31]), .B(A[31]), .Z(n323) );
  CND2X1 U422 ( .A(A[4]), .B(B[4]), .Z(n172) );
  CND2X1 U423 ( .A(A[10]), .B(B[10]), .Z(n141) );
  CND2X1 U424 ( .A(A[14]), .B(B[14]), .Z(n116) );
  CND2X1 U425 ( .A(A[12]), .B(B[12]), .Z(n128) );
  CND2X1 U426 ( .A(A[16]), .B(B[16]), .Z(n101) );
  CND2X1 U427 ( .A(A[2]), .B(B[2]), .Z(n181) );
  CND2X1 U428 ( .A(A[8]), .B(B[8]), .Z(n151) );
  CND2X1 U429 ( .A(A[18]), .B(B[18]), .Z(n91) );
  CND2X1 U430 ( .A(A[20]), .B(B[20]), .Z(n78) );
  CND2X1 U431 ( .A(A[22]), .B(B[22]), .Z(n70) );
  CND2X1 U432 ( .A(A[24]), .B(B[24]), .Z(n58) );
  CND2X1 U433 ( .A(A[26]), .B(B[26]), .Z(n48) );
  CND2X1 U434 ( .A(A[28]), .B(B[28]), .Z(n40) );
  CND2X1 U435 ( .A(A[21]), .B(B[21]), .Z(n75) );
  CND2X1 U436 ( .A(A[23]), .B(B[23]), .Z(n67) );
  CND2X1 U437 ( .A(A[27]), .B(B[27]), .Z(n43) );
  CND2X1 U438 ( .A(A[25]), .B(B[25]), .Z(n55) );
  COR2X1 U439 ( .A(A[26]), .B(B[26]), .Z(n324) );
  COR2X1 U440 ( .A(A[28]), .B(B[28]), .Z(n325) );
  CNR2X1 U441 ( .A(A[29]), .B(B[29]), .Z(n34) );
  CEOXL U442 ( .A(n187), .B(n30), .Z(n326) );
  CND2X1 U443 ( .A(A[29]), .B(B[29]), .Z(n35) );
  CIVX2 U444 ( .A(n101), .Z(n99) );
  CIVX2 U445 ( .A(n83), .Z(n81) );
  CIVX2 U446 ( .A(n48), .Z(n46) );
  CIVX2 U447 ( .A(n40), .Z(n38) );
  CIVX2 U448 ( .A(n184), .Z(n216) );
  CIVX2 U449 ( .A(n180), .Z(n215) );
  CIVX2 U450 ( .A(n177), .Z(n214) );
  CIVX2 U451 ( .A(n166), .Z(n212) );
  CIVX2 U452 ( .A(n161), .Z(n211) );
  CIVX2 U453 ( .A(n158), .Z(n210) );
  CIVX2 U454 ( .A(n150), .Z(n209) );
  CIVX2 U455 ( .A(n147), .Z(n208) );
  CIVX2 U456 ( .A(n135), .Z(n206) );
  CIVX2 U457 ( .A(n122), .Z(n204) );
  CIVX2 U458 ( .A(n110), .Z(n202) );
  CIVX2 U459 ( .A(n100), .Z(n98) );
  CIVX2 U460 ( .A(n95), .Z(n200) );
  CIVX2 U461 ( .A(n90), .Z(n199) );
  CIVX2 U462 ( .A(n87), .Z(n198) );
  CIVX2 U463 ( .A(n77), .Z(n197) );
  CIVX2 U464 ( .A(n74), .Z(n196) );
  CIVX2 U465 ( .A(n69), .Z(n195) );
  CIVX2 U466 ( .A(n66), .Z(n194) );
  CIVX2 U467 ( .A(n57), .Z(n193) );
  CIVX2 U468 ( .A(n54), .Z(n192) );
  CIVX2 U469 ( .A(n42), .Z(n190) );
  CIVX2 U470 ( .A(n34), .Z(n188) );
  CIVX2 U471 ( .A(n183), .Z(n182) );
  CIVX2 U472 ( .A(n174), .Z(n173) );
  CIVX2 U473 ( .A(n172), .Z(n170) );
  CIVX2 U474 ( .A(n171), .Z(n213) );
  CIVX2 U475 ( .A(n153), .Z(n152) );
  CIVX2 U476 ( .A(n146), .Z(n144) );
  CIVX2 U477 ( .A(n145), .Z(n143) );
  CIVX2 U478 ( .A(n141), .Z(n139) );
  CIVX2 U479 ( .A(n140), .Z(n207) );
  CIVX2 U480 ( .A(n130), .Z(n129) );
  CIVX2 U481 ( .A(n128), .Z(n126) );
  CIVX2 U482 ( .A(n127), .Z(n205) );
  CIVX2 U483 ( .A(n121), .Z(n119) );
  CIVX2 U484 ( .A(n120), .Z(n118) );
  CIVX2 U485 ( .A(n116), .Z(n114) );
  CIVX2 U486 ( .A(n115), .Z(n203) );
  CIVX2 U487 ( .A(n103), .Z(n102) );
endmodule


module calc_DW01_add_10 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n32, n33, n34, n35, n36, n38, n40, n41, n42, n43, n44, n46, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n187, n188, n190, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n326, n322, n323, n324, n325;

  CFA1X1 U3 ( .A(B[30]), .B(n33), .CI(A[30]), .CO(n32), .S(SUM[30]) );
  CAN2XL U252 ( .A(n322), .B(n187), .Z(SUM[0]) );
  CNIVX1 U253 ( .A(n326), .Z(SUM[1]) );
  COND1X2 U254 ( .A(n34), .B(n36), .C(n35), .Z(n33) );
  CANR1X1 U255 ( .A(n325), .B(n41), .C(n38), .Z(n36) );
  CANR1X1 U256 ( .A(n153), .B(n104), .C(n105), .Z(n103) );
  COND1X1 U257 ( .A(n154), .B(n174), .C(n155), .Z(n153) );
  CND2XL U258 ( .A(A[6]), .B(B[6]), .Z(n162) );
  COND1XL U259 ( .A(n42), .B(n44), .C(n43), .Z(n41) );
  CNR2XL U260 ( .A(n161), .B(n158), .Z(n156) );
  CANR1XL U261 ( .A(n52), .B(n61), .C(n53), .Z(n51) );
  COND1XL U262 ( .A(n187), .B(n184), .C(n185), .Z(n183) );
  CND2XL U263 ( .A(n216), .B(n185), .Z(n30) );
  CNR2X1 U264 ( .A(A[12]), .B(B[12]), .Z(n127) );
  CNR2XL U265 ( .A(n83), .B(n62), .Z(n60) );
  CIVX1 U266 ( .A(n80), .Z(n79) );
  CIVXL U267 ( .A(n84), .Z(n82) );
  COND1X1 U268 ( .A(n50), .B(n103), .C(n51), .Z(n49) );
  CND2XL U269 ( .A(n60), .B(n52), .Z(n50) );
  CND2XL U270 ( .A(n164), .B(n156), .Z(n154) );
  CNR2XL U271 ( .A(n127), .B(n122), .Z(n120) );
  CNR2XL U272 ( .A(n150), .B(n147), .Z(n145) );
  CNR2XL U273 ( .A(n90), .B(n87), .Z(n85) );
  CNR2XL U274 ( .A(n115), .B(n110), .Z(n108) );
  CNR2XL U275 ( .A(n140), .B(n135), .Z(n133) );
  CNR2XL U276 ( .A(n100), .B(n95), .Z(n93) );
  CEOXL U277 ( .A(n2), .B(n36), .Z(SUM[29]) );
  CND2XL U278 ( .A(n209), .B(n151), .Z(n23) );
  CND2XL U279 ( .A(n205), .B(n128), .Z(n19) );
  CND2XL U280 ( .A(n199), .B(n91), .Z(n13) );
  CND2XL U281 ( .A(n195), .B(n70), .Z(n9) );
  CEOXL U282 ( .A(n9), .B(n71), .Z(SUM[22]) );
  CEOXL U283 ( .A(n4), .B(n44), .Z(SUM[27]) );
  CND2XL U284 ( .A(n194), .B(n67), .Z(n8) );
  CND2XL U285 ( .A(n207), .B(n141), .Z(n21) );
  CND2XL U286 ( .A(n203), .B(n116), .Z(n17) );
  CND2XL U287 ( .A(n98), .B(n101), .Z(n15) );
  CND2XL U288 ( .A(n197), .B(n78), .Z(n11) );
  CND2XL U289 ( .A(n196), .B(n75), .Z(n10) );
  CEOXL U290 ( .A(n187), .B(n30), .Z(n326) );
  CND2XL U291 ( .A(n215), .B(n181), .Z(n29) );
  CND2XL U292 ( .A(n213), .B(n172), .Z(n27) );
  CNR2XL U293 ( .A(A[8]), .B(B[8]), .Z(n150) );
  CNR2XL U294 ( .A(A[16]), .B(B[16]), .Z(n100) );
  CND2XL U295 ( .A(A[1]), .B(B[1]), .Z(n185) );
  CND2XL U296 ( .A(A[3]), .B(B[3]), .Z(n178) );
  CND2XL U297 ( .A(A[9]), .B(B[9]), .Z(n148) );
  CND2XL U298 ( .A(A[13]), .B(B[13]), .Z(n123) );
  CND2XL U299 ( .A(A[7]), .B(B[7]), .Z(n159) );
  CND2XL U300 ( .A(A[5]), .B(B[5]), .Z(n167) );
  CND2XL U301 ( .A(A[11]), .B(B[11]), .Z(n136) );
  CND2XL U302 ( .A(A[15]), .B(B[15]), .Z(n111) );
  CND2XL U303 ( .A(A[19]), .B(B[19]), .Z(n88) );
  CND2XL U304 ( .A(A[17]), .B(B[17]), .Z(n96) );
  COR2XL U305 ( .A(A[0]), .B(B[0]), .Z(n322) );
  CANR1XL U306 ( .A(n164), .B(n173), .C(n165), .Z(n163) );
  CANR1XL U307 ( .A(n93), .B(n102), .C(n94), .Z(n92) );
  CANR1XL U308 ( .A(n72), .B(n79), .C(n73), .Z(n71) );
  CANR1XL U309 ( .A(n60), .B(n102), .C(n61), .Z(n59) );
  COND1XL U310 ( .A(n143), .B(n152), .C(n144), .Z(n142) );
  COND1XL U311 ( .A(n118), .B(n129), .C(n119), .Z(n117) );
  CNR2X1 U312 ( .A(n131), .B(n106), .Z(n104) );
  COND1XL U313 ( .A(n106), .B(n132), .C(n107), .Z(n105) );
  CND2X1 U314 ( .A(n120), .B(n108), .Z(n106) );
  CANR1XL U315 ( .A(n81), .B(n102), .C(n82), .Z(n80) );
  COND1XL U316 ( .A(n131), .B(n152), .C(n132), .Z(n130) );
  CND2X1 U317 ( .A(n93), .B(n85), .Z(n83) );
  CND2X1 U318 ( .A(n72), .B(n64), .Z(n62) );
  CND2X1 U319 ( .A(n145), .B(n133), .Z(n131) );
  CANR1XL U320 ( .A(n324), .B(n49), .C(n46), .Z(n44) );
  CNR2X1 U321 ( .A(n57), .B(n54), .Z(n52) );
  CENX1 U322 ( .A(n160), .B(n24), .Z(SUM[7]) );
  CND2X1 U323 ( .A(n210), .B(n159), .Z(n24) );
  COND1XL U324 ( .A(n161), .B(n163), .C(n162), .Z(n160) );
  CENX1 U325 ( .A(n68), .B(n8), .Z(SUM[23]) );
  COND1XL U326 ( .A(n69), .B(n71), .C(n70), .Z(n68) );
  CANR1XL U327 ( .A(n94), .B(n85), .C(n86), .Z(n84) );
  COND1XL U328 ( .A(n91), .B(n87), .C(n88), .Z(n86) );
  CANR1XL U329 ( .A(n183), .B(n175), .C(n176), .Z(n174) );
  CNR2X1 U330 ( .A(n180), .B(n177), .Z(n175) );
  COND1XL U331 ( .A(n181), .B(n177), .C(n178), .Z(n176) );
  CANR1XL U332 ( .A(n165), .B(n156), .C(n157), .Z(n155) );
  COND1XL U333 ( .A(n151), .B(n147), .C(n148), .Z(n146) );
  COND1XL U334 ( .A(n128), .B(n122), .C(n123), .Z(n121) );
  CANR1XL U335 ( .A(n146), .B(n133), .C(n134), .Z(n132) );
  COND1XL U336 ( .A(n141), .B(n135), .C(n136), .Z(n134) );
  COND1XL U337 ( .A(n172), .B(n166), .C(n167), .Z(n165) );
  COND1XL U338 ( .A(n101), .B(n95), .C(n96), .Z(n94) );
  COND1XL U339 ( .A(n78), .B(n74), .C(n75), .Z(n73) );
  COND1XL U340 ( .A(n62), .B(n84), .C(n63), .Z(n61) );
  CANR1XL U341 ( .A(n73), .B(n64), .C(n65), .Z(n63) );
  COND1XL U342 ( .A(n70), .B(n66), .C(n67), .Z(n65) );
  CANR1XL U343 ( .A(n121), .B(n108), .C(n109), .Z(n107) );
  COND1XL U344 ( .A(n116), .B(n110), .C(n111), .Z(n109) );
  CNR2X1 U345 ( .A(n69), .B(n66), .Z(n64) );
  CENX1 U346 ( .A(n149), .B(n22), .Z(SUM[9]) );
  CND2X1 U347 ( .A(n208), .B(n148), .Z(n22) );
  COND1XL U348 ( .A(n150), .B(n152), .C(n151), .Z(n149) );
  CENX1 U349 ( .A(n142), .B(n21), .Z(SUM[10]) );
  CENX1 U350 ( .A(n117), .B(n17), .Z(SUM[14]) );
  CENX1 U351 ( .A(n102), .B(n15), .Z(SUM[16]) );
  CENX1 U352 ( .A(n89), .B(n12), .Z(SUM[19]) );
  CND2X1 U353 ( .A(n198), .B(n88), .Z(n12) );
  COND1XL U354 ( .A(n90), .B(n92), .C(n91), .Z(n89) );
  CENX1 U355 ( .A(n79), .B(n11), .Z(SUM[20]) );
  CENX1 U356 ( .A(n76), .B(n10), .Z(SUM[21]) );
  COND1XL U357 ( .A(n77), .B(n80), .C(n78), .Z(n76) );
  CENX1 U358 ( .A(n56), .B(n6), .Z(SUM[25]) );
  CND2X1 U359 ( .A(n192), .B(n55), .Z(n6) );
  COND1XL U360 ( .A(n57), .B(n59), .C(n58), .Z(n56) );
  CENX1 U361 ( .A(n49), .B(n5), .Z(SUM[26]) );
  CND2X1 U362 ( .A(n324), .B(n48), .Z(n5) );
  CENX1 U363 ( .A(n41), .B(n3), .Z(SUM[28]) );
  CND2X1 U364 ( .A(n325), .B(n40), .Z(n3) );
  COND1XL U365 ( .A(n162), .B(n158), .C(n159), .Z(n157) );
  COND1XL U366 ( .A(n58), .B(n54), .C(n55), .Z(n53) );
  CNR2X1 U367 ( .A(n171), .B(n166), .Z(n164) );
  CNR2X1 U368 ( .A(n77), .B(n74), .Z(n72) );
  CEOX1 U369 ( .A(n20), .B(n137), .Z(SUM[11]) );
  CND2X1 U370 ( .A(n206), .B(n136), .Z(n20) );
  CANR1XL U371 ( .A(n207), .B(n142), .C(n139), .Z(n137) );
  CEOX1 U372 ( .A(n19), .B(n129), .Z(SUM[12]) );
  CEOX1 U373 ( .A(n18), .B(n124), .Z(SUM[13]) );
  CND2X1 U374 ( .A(n204), .B(n123), .Z(n18) );
  CANR1XL U375 ( .A(n205), .B(n130), .C(n126), .Z(n124) );
  CEOX1 U376 ( .A(n16), .B(n112), .Z(SUM[15]) );
  CND2X1 U377 ( .A(n202), .B(n111), .Z(n16) );
  CANR1XL U378 ( .A(n203), .B(n117), .C(n114), .Z(n112) );
  CEOX1 U379 ( .A(n14), .B(n97), .Z(SUM[17]) );
  CND2X1 U380 ( .A(n200), .B(n96), .Z(n14) );
  CANR1XL U381 ( .A(n98), .B(n102), .C(n99), .Z(n97) );
  CEOX1 U382 ( .A(n13), .B(n92), .Z(SUM[18]) );
  CEOX1 U383 ( .A(n7), .B(n59), .Z(SUM[24]) );
  CND2X1 U384 ( .A(n193), .B(n58), .Z(n7) );
  CND2X1 U385 ( .A(n190), .B(n43), .Z(n4) );
  CND2X1 U386 ( .A(n188), .B(n35), .Z(n2) );
  CEOX1 U387 ( .A(n26), .B(n168), .Z(SUM[5]) );
  CND2X1 U388 ( .A(n212), .B(n167), .Z(n26) );
  CANR1XL U389 ( .A(n213), .B(n173), .C(n170), .Z(n168) );
  CENX1 U390 ( .A(n179), .B(n28), .Z(SUM[3]) );
  CND2X1 U391 ( .A(n214), .B(n178), .Z(n28) );
  COND1XL U392 ( .A(n180), .B(n182), .C(n181), .Z(n179) );
  CENX1 U393 ( .A(n173), .B(n27), .Z(SUM[4]) );
  CEOX1 U394 ( .A(n29), .B(n182), .Z(SUM[2]) );
  CEOX1 U395 ( .A(n25), .B(n163), .Z(SUM[6]) );
  CND2X1 U396 ( .A(n211), .B(n162), .Z(n25) );
  CEOX1 U397 ( .A(n23), .B(n152), .Z(SUM[8]) );
  CNR2X1 U398 ( .A(A[5]), .B(B[5]), .Z(n166) );
  CNR2X1 U399 ( .A(A[17]), .B(B[17]), .Z(n95) );
  CNR2X1 U400 ( .A(A[19]), .B(B[19]), .Z(n87) );
  CNR2X1 U401 ( .A(A[21]), .B(B[21]), .Z(n74) );
  CNR2X1 U402 ( .A(A[23]), .B(B[23]), .Z(n66) );
  CNR2X1 U403 ( .A(A[9]), .B(B[9]), .Z(n147) );
  CNR2X1 U404 ( .A(A[3]), .B(B[3]), .Z(n177) );
  CNR2X1 U405 ( .A(A[11]), .B(B[11]), .Z(n135) );
  CNR2X1 U406 ( .A(A[15]), .B(B[15]), .Z(n110) );
  CNR2X1 U407 ( .A(A[13]), .B(B[13]), .Z(n122) );
  CNR2X1 U408 ( .A(A[7]), .B(B[7]), .Z(n158) );
  CNR2X1 U409 ( .A(A[25]), .B(B[25]), .Z(n54) );
  CNR2X1 U410 ( .A(A[2]), .B(B[2]), .Z(n180) );
  CNR2X1 U411 ( .A(A[6]), .B(B[6]), .Z(n161) );
  CNR2X1 U412 ( .A(A[18]), .B(B[18]), .Z(n90) );
  CNR2X1 U413 ( .A(A[20]), .B(B[20]), .Z(n77) );
  CNR2X1 U414 ( .A(A[22]), .B(B[22]), .Z(n69) );
  CNR2X1 U415 ( .A(A[24]), .B(B[24]), .Z(n57) );
  CNR2X1 U416 ( .A(A[14]), .B(B[14]), .Z(n115) );
  CNR2X1 U417 ( .A(A[10]), .B(B[10]), .Z(n140) );
  CNR2X1 U418 ( .A(A[4]), .B(B[4]), .Z(n171) );
  CND2X1 U419 ( .A(A[0]), .B(B[0]), .Z(n187) );
  CNR2X1 U420 ( .A(A[27]), .B(B[27]), .Z(n42) );
  CNR2X1 U421 ( .A(A[1]), .B(B[1]), .Z(n184) );
  CENX1 U422 ( .A(n323), .B(n32), .Z(SUM[31]) );
  CENX1 U423 ( .A(B[31]), .B(A[31]), .Z(n323) );
  CND2X1 U424 ( .A(A[4]), .B(B[4]), .Z(n172) );
  CND2X1 U425 ( .A(A[10]), .B(B[10]), .Z(n141) );
  CND2X1 U426 ( .A(A[14]), .B(B[14]), .Z(n116) );
  CND2X1 U427 ( .A(A[12]), .B(B[12]), .Z(n128) );
  CND2X1 U428 ( .A(A[16]), .B(B[16]), .Z(n101) );
  CND2X1 U429 ( .A(A[2]), .B(B[2]), .Z(n181) );
  CND2X1 U430 ( .A(A[8]), .B(B[8]), .Z(n151) );
  CND2X1 U431 ( .A(A[18]), .B(B[18]), .Z(n91) );
  CND2X1 U432 ( .A(A[20]), .B(B[20]), .Z(n78) );
  CND2X1 U433 ( .A(A[22]), .B(B[22]), .Z(n70) );
  CND2X1 U434 ( .A(A[24]), .B(B[24]), .Z(n58) );
  CND2X1 U435 ( .A(A[26]), .B(B[26]), .Z(n48) );
  CND2X1 U436 ( .A(A[28]), .B(B[28]), .Z(n40) );
  CND2X1 U437 ( .A(A[21]), .B(B[21]), .Z(n75) );
  CND2X1 U438 ( .A(A[23]), .B(B[23]), .Z(n67) );
  CND2X1 U439 ( .A(A[27]), .B(B[27]), .Z(n43) );
  CND2X1 U440 ( .A(A[25]), .B(B[25]), .Z(n55) );
  COR2X1 U441 ( .A(A[26]), .B(B[26]), .Z(n324) );
  COR2X1 U442 ( .A(A[28]), .B(B[28]), .Z(n325) );
  CNR2X1 U443 ( .A(A[29]), .B(B[29]), .Z(n34) );
  CND2X1 U444 ( .A(A[29]), .B(B[29]), .Z(n35) );
  CIVX2 U445 ( .A(n101), .Z(n99) );
  CIVX2 U446 ( .A(n83), .Z(n81) );
  CIVX2 U447 ( .A(n48), .Z(n46) );
  CIVX2 U448 ( .A(n40), .Z(n38) );
  CIVX2 U449 ( .A(n184), .Z(n216) );
  CIVX2 U450 ( .A(n180), .Z(n215) );
  CIVX2 U451 ( .A(n177), .Z(n214) );
  CIVX2 U452 ( .A(n166), .Z(n212) );
  CIVX2 U453 ( .A(n161), .Z(n211) );
  CIVX2 U454 ( .A(n158), .Z(n210) );
  CIVX2 U455 ( .A(n150), .Z(n209) );
  CIVX2 U456 ( .A(n147), .Z(n208) );
  CIVX2 U457 ( .A(n135), .Z(n206) );
  CIVX2 U458 ( .A(n122), .Z(n204) );
  CIVX2 U459 ( .A(n110), .Z(n202) );
  CIVX2 U460 ( .A(n100), .Z(n98) );
  CIVX2 U461 ( .A(n95), .Z(n200) );
  CIVX2 U462 ( .A(n90), .Z(n199) );
  CIVX2 U463 ( .A(n87), .Z(n198) );
  CIVX2 U464 ( .A(n77), .Z(n197) );
  CIVX2 U465 ( .A(n74), .Z(n196) );
  CIVX2 U466 ( .A(n69), .Z(n195) );
  CIVX2 U467 ( .A(n66), .Z(n194) );
  CIVX2 U468 ( .A(n57), .Z(n193) );
  CIVX2 U469 ( .A(n54), .Z(n192) );
  CIVX2 U470 ( .A(n42), .Z(n190) );
  CIVX2 U471 ( .A(n34), .Z(n188) );
  CIVX2 U472 ( .A(n183), .Z(n182) );
  CIVX2 U473 ( .A(n174), .Z(n173) );
  CIVX2 U474 ( .A(n172), .Z(n170) );
  CIVX2 U475 ( .A(n171), .Z(n213) );
  CIVX2 U476 ( .A(n153), .Z(n152) );
  CIVX2 U477 ( .A(n146), .Z(n144) );
  CIVX2 U478 ( .A(n145), .Z(n143) );
  CIVX2 U479 ( .A(n141), .Z(n139) );
  CIVX2 U480 ( .A(n140), .Z(n207) );
  CIVX2 U481 ( .A(n130), .Z(n129) );
  CIVX2 U482 ( .A(n128), .Z(n126) );
  CIVX2 U483 ( .A(n127), .Z(n205) );
  CIVX2 U484 ( .A(n121), .Z(n119) );
  CIVX2 U485 ( .A(n120), .Z(n118) );
  CIVX2 U486 ( .A(n116), .Z(n114) );
  CIVX2 U487 ( .A(n115), .Z(n203) );
  CIVX2 U488 ( .A(n103), .Z(n102) );
endmodule


module calc_DW01_add_11 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n38, n40, n41, n42, n43, n44, n46, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n190, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n324, n321, n322, n323;

  CFA1X1 U3 ( .A(B[30]), .B(n33), .CI(A[30]), .CO(n32), .S(SUM[30]) );
  CANR1X1 U252 ( .A(n323), .B(n41), .C(n38), .Z(n36) );
  COND1X1 U253 ( .A(n34), .B(n36), .C(n35), .Z(n33) );
  COND1X1 U254 ( .A(n154), .B(n174), .C(n155), .Z(n153) );
  CANR1X1 U255 ( .A(n183), .B(n175), .C(n176), .Z(n174) );
  CNIVX1 U256 ( .A(n324), .Z(SUM[1]) );
  CNR2X1 U257 ( .A(A[12]), .B(B[12]), .Z(n127) );
  CND2XL U258 ( .A(n120), .B(n108), .Z(n106) );
  CANR1XL U259 ( .A(n94), .B(n85), .C(n86), .Z(n84) );
  CND2XL U260 ( .A(n216), .B(n185), .Z(n30) );
  CNR2XL U261 ( .A(n83), .B(n62), .Z(n60) );
  CIVXL U262 ( .A(n80), .Z(n79) );
  CANR1X1 U263 ( .A(n153), .B(n104), .C(n105), .Z(n103) );
  COND1X1 U264 ( .A(n50), .B(n103), .C(n51), .Z(n49) );
  CND2XL U265 ( .A(n60), .B(n52), .Z(n50) );
  CANR1X1 U266 ( .A(n52), .B(n61), .C(n53), .Z(n51) );
  COND1X1 U267 ( .A(n42), .B(n44), .C(n43), .Z(n41) );
  CNR2XL U268 ( .A(n150), .B(n147), .Z(n145) );
  CNR2XL U269 ( .A(n127), .B(n122), .Z(n120) );
  CNR2XL U270 ( .A(n90), .B(n87), .Z(n85) );
  CNR2XL U271 ( .A(n140), .B(n135), .Z(n133) );
  CNR2XL U272 ( .A(n115), .B(n110), .Z(n108) );
  CNR2XL U273 ( .A(n69), .B(n66), .Z(n64) );
  CNR2XL U274 ( .A(n100), .B(n95), .Z(n93) );
  CNR2XL U275 ( .A(n171), .B(n166), .Z(n164) );
  CEOXL U276 ( .A(n2), .B(n36), .Z(SUM[29]) );
  CND2XL U277 ( .A(n211), .B(n162), .Z(n25) );
  CND2XL U278 ( .A(n209), .B(n151), .Z(n23) );
  CND2XL U279 ( .A(n205), .B(n128), .Z(n19) );
  CND2XL U280 ( .A(n199), .B(n91), .Z(n13) );
  CND2XL U281 ( .A(n195), .B(n70), .Z(n9) );
  CEOXL U282 ( .A(n9), .B(n71), .Z(SUM[22]) );
  CEOXL U283 ( .A(n4), .B(n44), .Z(SUM[27]) );
  CND2XL U284 ( .A(n207), .B(n141), .Z(n21) );
  CND2XL U285 ( .A(n203), .B(n116), .Z(n17) );
  CND2XL U286 ( .A(n98), .B(n101), .Z(n15) );
  CND2XL U287 ( .A(n197), .B(n78), .Z(n11) );
  CND2XL U288 ( .A(n196), .B(n75), .Z(n10) );
  CEOXL U289 ( .A(n187), .B(n30), .Z(n324) );
  CND2XL U290 ( .A(n215), .B(n181), .Z(n29) );
  CND2XL U291 ( .A(n213), .B(n172), .Z(n27) );
  CNR2XL U292 ( .A(A[8]), .B(B[8]), .Z(n150) );
  CNR2XL U293 ( .A(A[16]), .B(B[16]), .Z(n100) );
  CND2XL U294 ( .A(A[1]), .B(B[1]), .Z(n185) );
  CND2XL U295 ( .A(A[3]), .B(B[3]), .Z(n178) );
  CND2XL U296 ( .A(A[9]), .B(B[9]), .Z(n148) );
  CND2XL U297 ( .A(A[7]), .B(B[7]), .Z(n159) );
  CND2XL U298 ( .A(A[13]), .B(B[13]), .Z(n123) );
  CND2XL U299 ( .A(A[5]), .B(B[5]), .Z(n167) );
  CND2XL U300 ( .A(A[11]), .B(B[11]), .Z(n136) );
  CND2XL U301 ( .A(A[15]), .B(B[15]), .Z(n111) );
  CND2XL U302 ( .A(A[19]), .B(B[19]), .Z(n88) );
  CND2XL U303 ( .A(A[17]), .B(B[17]), .Z(n96) );
  CND2XL U304 ( .A(A[23]), .B(B[23]), .Z(n67) );
  CND2XL U305 ( .A(A[25]), .B(B[25]), .Z(n55) );
  CND2IXL U306 ( .B(n186), .A(n187), .Z(n31) );
  CNR2XL U307 ( .A(A[0]), .B(B[0]), .Z(n186) );
  CANR1XL U308 ( .A(n164), .B(n173), .C(n165), .Z(n163) );
  CANR1XL U309 ( .A(n93), .B(n102), .C(n94), .Z(n92) );
  CANR1XL U310 ( .A(n72), .B(n79), .C(n73), .Z(n71) );
  CANR1XL U311 ( .A(n60), .B(n102), .C(n61), .Z(n59) );
  COND1XL U312 ( .A(n143), .B(n152), .C(n144), .Z(n142) );
  COND1XL U313 ( .A(n118), .B(n129), .C(n119), .Z(n117) );
  CNR2X1 U314 ( .A(n131), .B(n106), .Z(n104) );
  COND1XL U315 ( .A(n106), .B(n132), .C(n107), .Z(n105) );
  CANR1XL U316 ( .A(n81), .B(n102), .C(n82), .Z(n80) );
  COND1XL U317 ( .A(n131), .B(n152), .C(n132), .Z(n130) );
  CND2X1 U318 ( .A(n93), .B(n85), .Z(n83) );
  CND2X1 U319 ( .A(n72), .B(n64), .Z(n62) );
  CND2X1 U320 ( .A(n145), .B(n133), .Z(n131) );
  CANR1XL U321 ( .A(n322), .B(n49), .C(n46), .Z(n44) );
  CNR2X1 U322 ( .A(n57), .B(n54), .Z(n52) );
  CENX1 U323 ( .A(n68), .B(n8), .Z(SUM[23]) );
  CND2X1 U324 ( .A(n194), .B(n67), .Z(n8) );
  COND1XL U325 ( .A(n69), .B(n71), .C(n70), .Z(n68) );
  COND1XL U326 ( .A(n91), .B(n87), .C(n88), .Z(n86) );
  CNR2X1 U327 ( .A(n180), .B(n177), .Z(n175) );
  COND1XL U328 ( .A(n181), .B(n177), .C(n178), .Z(n176) );
  COND1XL U329 ( .A(n128), .B(n122), .C(n123), .Z(n121) );
  CND2X1 U330 ( .A(n164), .B(n156), .Z(n154) );
  CANR1XL U331 ( .A(n165), .B(n156), .C(n157), .Z(n155) );
  CNR2X1 U332 ( .A(n161), .B(n158), .Z(n156) );
  COND1XL U333 ( .A(n187), .B(n184), .C(n185), .Z(n183) );
  COND1XL U334 ( .A(n151), .B(n147), .C(n148), .Z(n146) );
  CANR1XL U335 ( .A(n146), .B(n133), .C(n134), .Z(n132) );
  COND1XL U336 ( .A(n141), .B(n135), .C(n136), .Z(n134) );
  COND1XL U337 ( .A(n172), .B(n166), .C(n167), .Z(n165) );
  COND1XL U338 ( .A(n101), .B(n95), .C(n96), .Z(n94) );
  COND1XL U339 ( .A(n78), .B(n74), .C(n75), .Z(n73) );
  COND1XL U340 ( .A(n62), .B(n84), .C(n63), .Z(n61) );
  CANR1XL U341 ( .A(n73), .B(n64), .C(n65), .Z(n63) );
  COND1XL U342 ( .A(n70), .B(n66), .C(n67), .Z(n65) );
  CANR1XL U343 ( .A(n121), .B(n108), .C(n109), .Z(n107) );
  COND1XL U344 ( .A(n116), .B(n110), .C(n111), .Z(n109) );
  CENX1 U345 ( .A(n160), .B(n24), .Z(SUM[7]) );
  CND2X1 U346 ( .A(n210), .B(n159), .Z(n24) );
  COND1XL U347 ( .A(n161), .B(n163), .C(n162), .Z(n160) );
  CENX1 U348 ( .A(n149), .B(n22), .Z(SUM[9]) );
  CND2X1 U349 ( .A(n208), .B(n148), .Z(n22) );
  COND1XL U350 ( .A(n150), .B(n152), .C(n151), .Z(n149) );
  CENX1 U351 ( .A(n142), .B(n21), .Z(SUM[10]) );
  CENX1 U352 ( .A(n117), .B(n17), .Z(SUM[14]) );
  CENX1 U353 ( .A(n102), .B(n15), .Z(SUM[16]) );
  CENX1 U354 ( .A(n89), .B(n12), .Z(SUM[19]) );
  CND2X1 U355 ( .A(n198), .B(n88), .Z(n12) );
  COND1XL U356 ( .A(n90), .B(n92), .C(n91), .Z(n89) );
  CENX1 U357 ( .A(n79), .B(n11), .Z(SUM[20]) );
  CENX1 U358 ( .A(n76), .B(n10), .Z(SUM[21]) );
  COND1XL U359 ( .A(n77), .B(n80), .C(n78), .Z(n76) );
  CENX1 U360 ( .A(n56), .B(n6), .Z(SUM[25]) );
  CND2X1 U361 ( .A(n192), .B(n55), .Z(n6) );
  COND1XL U362 ( .A(n57), .B(n59), .C(n58), .Z(n56) );
  CENX1 U363 ( .A(n49), .B(n5), .Z(SUM[26]) );
  CND2X1 U364 ( .A(n322), .B(n48), .Z(n5) );
  CENX1 U365 ( .A(n41), .B(n3), .Z(SUM[28]) );
  CND2X1 U366 ( .A(n323), .B(n40), .Z(n3) );
  COND1XL U367 ( .A(n162), .B(n158), .C(n159), .Z(n157) );
  COND1XL U368 ( .A(n58), .B(n54), .C(n55), .Z(n53) );
  CNR2X1 U369 ( .A(n77), .B(n74), .Z(n72) );
  CEOX1 U370 ( .A(n20), .B(n137), .Z(SUM[11]) );
  CND2X1 U371 ( .A(n206), .B(n136), .Z(n20) );
  CANR1XL U372 ( .A(n207), .B(n142), .C(n139), .Z(n137) );
  CEOX1 U373 ( .A(n19), .B(n129), .Z(SUM[12]) );
  CEOX1 U374 ( .A(n18), .B(n124), .Z(SUM[13]) );
  CND2X1 U375 ( .A(n204), .B(n123), .Z(n18) );
  CANR1XL U376 ( .A(n205), .B(n130), .C(n126), .Z(n124) );
  CEOX1 U377 ( .A(n16), .B(n112), .Z(SUM[15]) );
  CND2X1 U378 ( .A(n202), .B(n111), .Z(n16) );
  CANR1XL U379 ( .A(n203), .B(n117), .C(n114), .Z(n112) );
  CEOX1 U380 ( .A(n14), .B(n97), .Z(SUM[17]) );
  CND2X1 U381 ( .A(n200), .B(n96), .Z(n14) );
  CANR1XL U382 ( .A(n98), .B(n102), .C(n99), .Z(n97) );
  CEOX1 U383 ( .A(n13), .B(n92), .Z(SUM[18]) );
  CEOX1 U384 ( .A(n7), .B(n59), .Z(SUM[24]) );
  CND2X1 U385 ( .A(n193), .B(n58), .Z(n7) );
  CND2X1 U386 ( .A(n190), .B(n43), .Z(n4) );
  CND2X1 U387 ( .A(n188), .B(n35), .Z(n2) );
  CEOX1 U388 ( .A(n26), .B(n168), .Z(SUM[5]) );
  CND2X1 U389 ( .A(n212), .B(n167), .Z(n26) );
  CANR1XL U390 ( .A(n213), .B(n173), .C(n170), .Z(n168) );
  CENX1 U391 ( .A(n179), .B(n28), .Z(SUM[3]) );
  CND2X1 U392 ( .A(n214), .B(n178), .Z(n28) );
  COND1XL U393 ( .A(n180), .B(n182), .C(n181), .Z(n179) );
  CENX1 U394 ( .A(n173), .B(n27), .Z(SUM[4]) );
  CEOX1 U395 ( .A(n29), .B(n182), .Z(SUM[2]) );
  CEOX1 U396 ( .A(n25), .B(n163), .Z(SUM[6]) );
  CEOX1 U397 ( .A(n23), .B(n152), .Z(SUM[8]) );
  CNR2X1 U398 ( .A(A[5]), .B(B[5]), .Z(n166) );
  CNR2X1 U399 ( .A(A[7]), .B(B[7]), .Z(n158) );
  CNR2X1 U400 ( .A(A[13]), .B(B[13]), .Z(n122) );
  CNR2X1 U401 ( .A(A[15]), .B(B[15]), .Z(n110) );
  CNR2X1 U402 ( .A(A[17]), .B(B[17]), .Z(n95) );
  CNR2X1 U403 ( .A(A[19]), .B(B[19]), .Z(n87) );
  CNR2X1 U404 ( .A(A[21]), .B(B[21]), .Z(n74) );
  CNR2X1 U405 ( .A(A[23]), .B(B[23]), .Z(n66) );
  CNR2X1 U406 ( .A(A[3]), .B(B[3]), .Z(n177) );
  CNR2X1 U407 ( .A(A[11]), .B(B[11]), .Z(n135) );
  CNR2X1 U408 ( .A(A[9]), .B(B[9]), .Z(n147) );
  CNR2X1 U409 ( .A(A[25]), .B(B[25]), .Z(n54) );
  CNR2X1 U410 ( .A(A[2]), .B(B[2]), .Z(n180) );
  CNR2X1 U411 ( .A(A[6]), .B(B[6]), .Z(n161) );
  CNR2X1 U412 ( .A(A[18]), .B(B[18]), .Z(n90) );
  CNR2X1 U413 ( .A(A[20]), .B(B[20]), .Z(n77) );
  CNR2X1 U414 ( .A(A[22]), .B(B[22]), .Z(n69) );
  CNR2X1 U415 ( .A(A[24]), .B(B[24]), .Z(n57) );
  CNR2X1 U416 ( .A(A[10]), .B(B[10]), .Z(n140) );
  CNR2X1 U417 ( .A(A[4]), .B(B[4]), .Z(n171) );
  CNR2X1 U418 ( .A(A[14]), .B(B[14]), .Z(n115) );
  CND2X1 U419 ( .A(A[0]), .B(B[0]), .Z(n187) );
  CNR2X1 U420 ( .A(A[27]), .B(B[27]), .Z(n42) );
  CNR2X1 U421 ( .A(A[1]), .B(B[1]), .Z(n184) );
  CENX1 U422 ( .A(n321), .B(n32), .Z(SUM[31]) );
  CENX1 U423 ( .A(B[31]), .B(A[31]), .Z(n321) );
  CND2X1 U424 ( .A(A[4]), .B(B[4]), .Z(n172) );
  CND2X1 U425 ( .A(A[10]), .B(B[10]), .Z(n141) );
  CND2X1 U426 ( .A(A[14]), .B(B[14]), .Z(n116) );
  CND2X1 U427 ( .A(A[12]), .B(B[12]), .Z(n128) );
  CND2X1 U428 ( .A(A[16]), .B(B[16]), .Z(n101) );
  CND2X1 U429 ( .A(A[2]), .B(B[2]), .Z(n181) );
  CND2X1 U430 ( .A(A[6]), .B(B[6]), .Z(n162) );
  CND2X1 U431 ( .A(A[8]), .B(B[8]), .Z(n151) );
  CND2X1 U432 ( .A(A[18]), .B(B[18]), .Z(n91) );
  CND2X1 U433 ( .A(A[20]), .B(B[20]), .Z(n78) );
  CND2X1 U434 ( .A(A[22]), .B(B[22]), .Z(n70) );
  CND2X1 U435 ( .A(A[24]), .B(B[24]), .Z(n58) );
  CND2X1 U436 ( .A(A[26]), .B(B[26]), .Z(n48) );
  CND2X1 U437 ( .A(A[28]), .B(B[28]), .Z(n40) );
  CND2X1 U438 ( .A(A[21]), .B(B[21]), .Z(n75) );
  CND2X1 U439 ( .A(A[27]), .B(B[27]), .Z(n43) );
  COR2X1 U440 ( .A(A[26]), .B(B[26]), .Z(n322) );
  COR2X1 U441 ( .A(A[28]), .B(B[28]), .Z(n323) );
  CNR2X1 U442 ( .A(A[29]), .B(B[29]), .Z(n34) );
  CND2X1 U443 ( .A(A[29]), .B(B[29]), .Z(n35) );
  CIVX2 U444 ( .A(n101), .Z(n99) );
  CIVX2 U445 ( .A(n84), .Z(n82) );
  CIVX2 U446 ( .A(n83), .Z(n81) );
  CIVX2 U447 ( .A(n48), .Z(n46) );
  CIVX2 U448 ( .A(n40), .Z(n38) );
  CIVX2 U449 ( .A(n184), .Z(n216) );
  CIVX2 U450 ( .A(n180), .Z(n215) );
  CIVX2 U451 ( .A(n177), .Z(n214) );
  CIVX2 U452 ( .A(n166), .Z(n212) );
  CIVX2 U453 ( .A(n161), .Z(n211) );
  CIVX2 U454 ( .A(n158), .Z(n210) );
  CIVX2 U455 ( .A(n150), .Z(n209) );
  CIVX2 U456 ( .A(n147), .Z(n208) );
  CIVX2 U457 ( .A(n135), .Z(n206) );
  CIVX2 U458 ( .A(n122), .Z(n204) );
  CIVX2 U459 ( .A(n110), .Z(n202) );
  CIVX2 U460 ( .A(n100), .Z(n98) );
  CIVX2 U461 ( .A(n95), .Z(n200) );
  CIVX2 U462 ( .A(n90), .Z(n199) );
  CIVX2 U463 ( .A(n87), .Z(n198) );
  CIVX2 U464 ( .A(n77), .Z(n197) );
  CIVX2 U465 ( .A(n74), .Z(n196) );
  CIVX2 U466 ( .A(n69), .Z(n195) );
  CIVX2 U467 ( .A(n66), .Z(n194) );
  CIVX2 U468 ( .A(n57), .Z(n193) );
  CIVX2 U469 ( .A(n54), .Z(n192) );
  CIVX2 U470 ( .A(n42), .Z(n190) );
  CIVX2 U471 ( .A(n34), .Z(n188) );
  CIVX2 U472 ( .A(n183), .Z(n182) );
  CIVX2 U473 ( .A(n174), .Z(n173) );
  CIVX2 U474 ( .A(n172), .Z(n170) );
  CIVX2 U475 ( .A(n171), .Z(n213) );
  CIVX2 U476 ( .A(n153), .Z(n152) );
  CIVX2 U477 ( .A(n146), .Z(n144) );
  CIVX2 U478 ( .A(n145), .Z(n143) );
  CIVX2 U479 ( .A(n141), .Z(n139) );
  CIVX2 U480 ( .A(n140), .Z(n207) );
  CIVX2 U481 ( .A(n130), .Z(n129) );
  CIVX2 U482 ( .A(n128), .Z(n126) );
  CIVX2 U483 ( .A(n127), .Z(n205) );
  CIVX2 U484 ( .A(n121), .Z(n119) );
  CIVX2 U485 ( .A(n120), .Z(n118) );
  CIVX2 U486 ( .A(n116), .Z(n114) );
  CIVX2 U487 ( .A(n115), .Z(n203) );
  CIVX2 U488 ( .A(n103), .Z(n102) );
  CIVX2 U489 ( .A(n31), .Z(SUM[0]) );
endmodule


module calc_DW_mult_tc_23 ( a, b, product, i_retiming_group_0_clk );
  input [32:0] a;
  input [32:0] b;
  output [65:0] product;
  input i_retiming_group_0_clk;
  wire   n3, n6, n9, n12, n18, n21, n27, n30, n33, n36, n39, n42, n44, n48,
         n50, n53, n55, n58, n61, n63, n66, n69, n71, n74, n77, n79, n84, n86,
         n89, n91, n93, n95, n97, n99, n100, n102, n104, n105, n107, n109,
         n110, n112, n113, n116, n120, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n157, n162, n164,
         n165, n166, n167, n171, n172, n179, n180, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n192, n194, n195, n196, n197, n201,
         n203, n204, n205, n206, n207, n208, n212, n214, n215, n216, n217,
         n219, n222, n223, n224, n225, n227, n229, n230, n231, n232, n233,
         n234, n235, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n250, n252, n253, n254, n255, n257, n260, n261,
         n262, n263, n265, n267, n268, n269, n270, n271, n272, n273, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n288, n289, n290, n292, n294, n295, n297, n299, n300, n301, n303,
         n305, n306, n307, n308, n309, n311, n313, n314, n315, n316, n317,
         n319, n321, n322, n323, n324, n325, n327, n329, n330, n332, n335,
         n336, n337, n338, n342, n344, n345, n346, n348, n350, n351, n353,
         n361, n364, n365, n366, n367, n368, n369, n370, n373, n375, n378,
         n379, n381, n382, n383, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n411, n412, n417, n418, n419, n421, n423,
         n424, n425, n426, n427, n428, n429, n430, n434, n435, n437, n438,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1407, n1408, n1409, n1410, n1411,
         n1412, n1415, n1416, n1417, n1418, n1420, n1421, n1432, n1435, n1436,
         n1438, n2259, n2258, n2257, net33082, net33080, net33480, net33482,
         net171503, net171634, net171635, net171637, net171639, net171643,
         net171708, net171723, net171725, net171738, net171752, net171759,
         net179371, net179544, net179680, net179686, net179834, net179913,
         net179912, net179947, net179954, net179996, net180018, net180017,
         net180016, net180095, net180094, net180107, net180106, net180105,
         net180475, net180482, net180480, net179493, net179380, n151, n1431,
         n1406, n115, n114, n1088, n1087, n1086, net182663, net182662,
         net184228, net182724, n420, net180013, net179971, net179515,
         net179430, net179197, net178620, n178, n175, n173, n160, n159, n158,
         n156, n154, n152, net179910, net179805, n464, n463, n462, n461, n439,
         n436, n422, n416, n415, n414, n413, n410, n409, n408, n407, n384,
         n380, n163, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1629, n1631, n1632, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256;
  assign n3 = a[1];
  assign n12 = a[3];
  assign n21 = a[5];
  assign n30 = a[7];
  assign n39 = a[9];
  assign n48 = a[11];
  assign n55 = a[13];
  assign n63 = a[15];
  assign n71 = a[17];
  assign n79 = a[19];
  assign n86 = a[21];
  assign n93 = a[23];
  assign n99 = a[25];
  assign n104 = a[27];
  assign n109 = a[29];
  assign n113 = a[32];
  assign n116 = b[0];
  assign n1382 = b[23];
  assign n1383 = b[22];
  assign n1384 = b[21];
  assign n1385 = b[20];
  assign n1386 = b[19];
  assign n1387 = b[18];
  assign n1388 = b[17];
  assign n1389 = b[16];
  assign n1390 = b[15];
  assign n1391 = b[14];
  assign n1392 = b[13];
  assign n1393 = b[12];
  assign n1394 = b[11];
  assign n1395 = b[10];
  assign n1396 = b[9];
  assign n1397 = b[8];
  assign n1398 = b[7];
  assign n1399 = b[6];
  assign n1400 = b[5];
  assign n1401 = b[4];
  assign n1402 = b[3];
  assign n1403 = b[2];
  assign n1404 = b[1];
  assign n2183 = i_retiming_group_0_clk;

  CEO3X2 U371 ( .A(n383), .B(n365), .C(n381), .Z(n364) );
  CEO3X2 U372 ( .A(n385), .B(n367), .C(n366), .Z(n365) );
  CEO3X2 U373 ( .A(n369), .B(n387), .C(n368), .Z(n366) );
  CEO3X2 U374 ( .A(n391), .B(n370), .C(n389), .Z(n367) );
  CEO3X2 U380 ( .A(n971), .B(n997), .C(n1025), .Z(n373) );
  CEO3X2 U382 ( .A(n2083), .B(n2064), .C(n2041), .Z(n375) );
  CFA1X1 U387 ( .A(n388), .B(n386), .CI(n411), .CO(n381), .S(n382) );
  CFA1X1 U389 ( .A(n417), .B(n392), .CI(n394), .CO(n385), .S(n386) );
  CFA1X1 U390 ( .A(n421), .B(n396), .CI(n419), .CO(n387), .S(n388) );
  CFA1X1 U391 ( .A(n402), .B(n2158), .CI(n2153), .CO(n389), .S(n390) );
  CFA1X1 U392 ( .A(n2154), .B(n404), .CI(n2156), .CO(n391), .S(n392) );
  CFA1X1 U394 ( .A(n2034), .B(n429), .CI(n2165), .CO(n395), .S(n396) );
  CFA1X1 U395 ( .A(n972), .B(n1056), .CI(n1026), .CO(n397), .S(n398) );
  CFA1X1 U397 ( .A(n2082), .B(n2042), .CI(n2085), .CO(n401), .S(n402) );
  CFA1X1 U398 ( .A(n2076), .B(n2057), .CI(n2061), .CO(n403), .S(n404) );
  CFA1X1 U402 ( .A(n443), .B(n441), .CI(n418), .CO(n411), .S(n412) );
  CFA1X1 U408 ( .A(n999), .B(n434), .CI(n1027), .CO(n423), .S(n424) );
  CFA1X1 U410 ( .A(n859), .B(n949), .CI(n889), .CO(n427), .S(n428) );
  CFA1X1 U411 ( .A(n2075), .B(n2043), .CI(n2081), .CO(n429), .S(n430) );
  CFA1X1 U415 ( .A(n444), .B(n442), .CI(n465), .CO(n437), .S(n438) );
  CFA1X1 U418 ( .A(n2151), .B(n473), .CI(n475), .CO(n443), .S(n444) );
  CFA1X1 U422 ( .A(n974), .B(n1058), .CI(n1000), .CO(n451), .S(n452) );
  CFA1X1 U423 ( .A(n890), .B(n1028), .CI(n950), .CO(n453), .S(n454) );
  CFA1X1 U431 ( .A(n482), .B(n499), .CI(n2148), .CO(n469), .S(n470) );
  CFA1X1 U433 ( .A(n2144), .B(n505), .CI(n2146), .CO(n473), .S(n474) );
  CFA1X1 U435 ( .A(n975), .B(n1059), .CI(n1029), .CO(n477), .S(n478) );
  CHA1X1 U439 ( .A(n849), .B(n875), .CO(n485), .S(n486) );
  CFA1X1 U447 ( .A(n976), .B(n533), .CI(n1002), .CO(n501), .S(n502) );
  CFA1X1 U448 ( .A(n952), .B(n1060), .CI(n1030), .CO(n503), .S(n504) );
  CFA1X1 U453 ( .A(n541), .B(n539), .CI(n518), .CO(n513), .S(n514) );
  CFA1X1 U459 ( .A(n977), .B(n1031), .CI(n1003), .CO(n525), .S(n526) );
  CHA1X1 U463 ( .A(n851), .B(n893), .CO(n533), .S(n534) );
  CFA1X1 U465 ( .A(n563), .B(n542), .CI(n561), .CO(n537), .S(n538) );
  CFA1X1 U467 ( .A(n2129), .B(n2136), .CI(n567), .CO(n541), .S(n542) );
  CFA1X1 U468 ( .A(n2132), .B(n2135), .CI(n2134), .CO(n543), .S(n544) );
  CFA1X1 U470 ( .A(n1004), .B(n575), .CI(n577), .CO(n547), .S(n548) );
  CFA1X1 U471 ( .A(n1062), .B(n978), .CI(n1032), .CO(n549), .S(n550) );
  CFA1X1 U474 ( .A(n834), .B(n864), .CI(n852), .CO(n555), .S(n556) );
  CFA1X1 U475 ( .A(n562), .B(n560), .CI(n581), .CO(n557), .S(n558) );
  CFA1X1 U477 ( .A(n587), .B(n585), .CI(n568), .CO(n561), .S(n562) );
  CFA1X1 U480 ( .A(n2118), .B(n2122), .CI(n2120), .CO(n567), .S(n568) );
  CFA1X1 U486 ( .A(n584), .B(n582), .CI(n601), .CO(n579), .S(n580) );
  CFA1X1 U487 ( .A(n588), .B(n603), .CI(n586), .CO(n581), .S(n582) );
  CFA1X1 U489 ( .A(n2121), .B(n2116), .CI(n2123), .CO(n585), .S(n586) );
  CFA1X1 U490 ( .A(n2160), .B(n2119), .CI(n2117), .CO(n587), .S(n588) );
  CFA1X1 U492 ( .A(n980), .B(n1034), .CI(n1006), .CO(n591), .S(n592) );
  CFA1X1 U493 ( .A(n914), .B(n1064), .CI(n934), .CO(n593), .S(n594) );
  CFA1X1 U496 ( .A(n604), .B(n602), .CI(n621), .CO(n599), .S(n600) );
  CFA1X1 U497 ( .A(n608), .B(n623), .CI(n606), .CO(n601), .S(n602) );
  CFA1X1 U498 ( .A(n2108), .B(n2110), .CI(n2115), .CO(n603), .S(n604) );
  CFA1X1 U499 ( .A(n2106), .B(n2169), .CI(n2113), .CO(n605), .S(n606) );
  CFA1X1 U500 ( .A(n2103), .B(n2111), .CI(n2104), .CO(n607), .S(n608) );
  CFA1X1 U503 ( .A(n935), .B(n1065), .CI(n915), .CO(n613), .S(n614) );
  CFA1X1 U504 ( .A(n881), .B(n957), .CI(n804), .CO(n615), .S(n616) );
  CFA1X1 U506 ( .A(n624), .B(n622), .CI(n639), .CO(n619), .S(n620) );
  CFA1X1 U507 ( .A(n2107), .B(n2102), .CI(n2109), .CO(n621), .S(n622) );
  CFA1X1 U508 ( .A(n2105), .B(n643), .CI(n2100), .CO(n623), .S(n624) );
  CFA1X1 U511 ( .A(n958), .B(n653), .CI(n982), .CO(n629), .S(n630) );
  CFA1X1 U512 ( .A(n1066), .B(n936), .CI(n1008), .CO(n631), .S(n632) );
  CFA1X1 U514 ( .A(n882), .B(n868), .CI(n856), .CO(n635), .S(n636) );
  CFA1X1 U515 ( .A(n2101), .B(n640), .CI(n2097), .CO(n637), .S(n638) );
  CFA1X1 U516 ( .A(n2099), .B(n2095), .CI(n644), .CO(n639), .S(n640) );
  CFA1X1 U517 ( .A(n648), .B(n661), .CI(n663), .CO(n641), .S(n642) );
  CFA1X1 U518 ( .A(n2093), .B(n2039), .CI(n2098), .CO(n643), .S(n644) );
  CFA1X1 U519 ( .A(n654), .B(n667), .CI(n669), .CO(n645), .S(n646) );
  CFA1X1 U520 ( .A(n959), .B(n1037), .CI(n983), .CO(n647), .S(n648) );
  CHA1X1 U523 ( .A(n883), .B(n917), .CO(n653), .S(n654) );
  CFA1X1 U524 ( .A(n2094), .B(n2096), .CI(n2090), .CO(n655), .S(n656) );
  CFA1X1 U526 ( .A(n666), .B(n677), .CI(n679), .CO(n659), .S(n660) );
  CFA1X1 U528 ( .A(n984), .B(n683), .CI(n685), .CO(n663), .S(n664) );
  CFA1X1 U529 ( .A(n938), .B(n1038), .CI(n1010), .CO(n665), .S(n666) );
  CFA1X1 U530 ( .A(n918), .B(n1068), .CI(n960), .CO(n667), .S(n668) );
  CFA1X1 U536 ( .A(n1011), .B(n686), .CI(n1039), .CO(n679), .S(n680) );
  CFA1X1 U537 ( .A(n919), .B(n885), .CI(n985), .CO(n681), .S(n682) );
  CFA1X1 U540 ( .A(n692), .B(n690), .CI(n703), .CO(n687), .S(n688) );
  CFA1X1 U541 ( .A(n707), .B(n694), .CI(n705), .CO(n689), .S(n690) );
  CFA1X1 U543 ( .A(n713), .B(n709), .CI(n711), .CO(n693), .S(n694) );
  CFA1X1 U544 ( .A(n962), .B(n1040), .CI(n986), .CO(n695), .S(n696) );
  CFA1X1 U545 ( .A(n1609), .B(n1070), .CI(n1012), .CO(n697), .S(n698) );
  CFA1X1 U546 ( .A(n886), .B(n920), .CI(n902), .CO(n699), .S(n700) );
  CFA1X1 U550 ( .A(n1013), .B(n714), .CI(n725), .CO(n707), .S(n708) );
  CFA1X1 U554 ( .A(n720), .B(n718), .CI(n729), .CO(n715), .S(n716) );
  CFA1X1 U555 ( .A(n724), .B(n731), .CI(n722), .CO(n717), .S(n718) );
  CFA1X1 U556 ( .A(n735), .B(n726), .CI(n733), .CO(n719), .S(n720) );
  CFA1X1 U557 ( .A(n988), .B(n737), .CI(n1014), .CO(n721), .S(n722) );
  CFA1X1 U560 ( .A(n732), .B(n730), .CI(n741), .CO(n727), .S(n728) );
  CFA1X1 U561 ( .A(n736), .B(n743), .CI(n734), .CO(n729), .S(n730) );
  CFA1X1 U562 ( .A(n738), .B(n745), .CI(n747), .CO(n731), .S(n732) );
  CFA1X1 U563 ( .A(n989), .B(n923), .CI(n1043), .CO(n733), .S(n734) );
  CHA1X1 U565 ( .A(n808), .B(n965), .CO(n737), .S(n738) );
  CFA1X1 U568 ( .A(n1016), .B(n755), .CI(n757), .CO(n743), .S(n744) );
  CFA1X1 U569 ( .A(n990), .B(n1074), .CI(n1044), .CO(n745), .S(n746) );
  CFA1X1 U570 ( .A(n924), .B(n966), .CI(n944), .CO(n747), .S(n748) );
  CFA1X1 U571 ( .A(n754), .B(n752), .CI(n761), .CO(n749), .S(n750) );
  CFA1X1 U572 ( .A(n765), .B(n756), .CI(n763), .CO(n751), .S(n752) );
  CFA1X1 U576 ( .A(n764), .B(n762), .CI(n769), .CO(n759), .S(n760) );
  CFA1X1 U577 ( .A(n773), .B(n766), .CI(n771), .CO(n761), .S(n762) );
  CFA1X1 U580 ( .A(n777), .B(n770), .CI(n772), .CO(n767), .S(n768) );
  CFA1X1 U581 ( .A(n1019), .B(n779), .CI(n774), .CO(n769), .S(n770) );
  CFA1X1 U582 ( .A(n969), .B(n1047), .CI(n993), .CO(n771), .S(n772) );
  CFA1X1 U584 ( .A(n783), .B(n778), .CI(n780), .CO(n775), .S(n776) );
  CFA1X1 U585 ( .A(n1048), .B(n785), .CI(n1078), .CO(n777), .S(n778) );
  CFA1X1 U587 ( .A(n786), .B(n784), .CI(n789), .CO(n781), .S(n782) );
  CFA1X1 U590 ( .A(n1080), .B(n790), .CI(n793), .CO(n787), .S(n788) );
  CFA1X1 U591 ( .A(n996), .B(n1050), .CI(n1022), .CO(n789), .S(n790) );
  CFA1X1 U592 ( .A(n1051), .B(n794), .CI(n1081), .CO(n791), .S(n792) );
  CHA1X1 U593 ( .A(n812), .B(n1023), .CO(n793), .S(n794) );
  CFA1X1 U594 ( .A(n1024), .B(n1082), .CI(n1052), .CO(n795), .S(n796) );
  CHA1X1 U595 ( .A(n813), .B(n1083), .CO(n797), .S(n798) );
  COND2X1 U646 ( .A(n97), .B(n1112), .C(n95), .D(n1111), .Z(n836) );
  COND2X1 U675 ( .A(n1964), .B(n1130), .C(n89), .D(n1692), .Z(n853) );
  COND2X1 U704 ( .A(n1905), .B(n1146), .C(n1865), .D(n1145), .Z(n868) );
  COND2X1 U722 ( .A(n1970), .B(n1438), .C(n74), .D(n1165), .Z(n806) );
  CND2IX1 U835 ( .B(net33082), .A(n2255), .Z(n1205) );
  COND2X1 U903 ( .A(n44), .B(n1250), .C(n1249), .D(n42), .Z(n967) );
  COND2X1 U905 ( .A(n1252), .B(n44), .C(n42), .D(n1251), .Z(n969) );
  COND2X1 U951 ( .A(n36), .B(n1273), .C(n1272), .D(n33), .Z(n989) );
  COND2X1 U955 ( .A(n36), .B(n1277), .C(n1276), .D(n33), .Z(n993) );
  COND2X1 U956 ( .A(n36), .B(n1278), .C(n1277), .D(n33), .Z(n994) );
  COND2X1 U1005 ( .A(n27), .B(n1300), .C(n1299), .D(n2009), .Z(n1015) );
  COND2X1 U1064 ( .A(n18), .B(n1330), .C(n1329), .D(n2185), .Z(n1044) );
  COND2X1 U1072 ( .A(n18), .B(n1338), .C(n1337), .D(n2185), .Z(n1052) );
  COND2X1 U1107 ( .A(n9), .B(n1342), .C(n6), .D(n1341), .Z(n1055) );
  COND2X1 U1108 ( .A(n9), .B(n1343), .C(n6), .D(n1342), .Z(n1056) );
  COND2X1 U1109 ( .A(n9), .B(n1344), .C(n6), .D(n1343), .Z(n1057) );
  COND2X1 U1110 ( .A(n9), .B(n1345), .C(n6), .D(n1344), .Z(n1058) );
  COND2X1 U1111 ( .A(n9), .B(n1346), .C(n6), .D(n1345), .Z(n1059) );
  COND2X1 U1112 ( .A(n9), .B(n1347), .C(n6), .D(n1346), .Z(n1060) );
  COND2X1 U1114 ( .A(n9), .B(n1349), .C(n6), .D(n1348), .Z(n1062) );
  COND2X1 U1116 ( .A(n9), .B(n1351), .C(n6), .D(n1350), .Z(n1064) );
  COND2X1 U1117 ( .A(n9), .B(n1352), .C(n6), .D(n1351), .Z(n1065) );
  COND2X1 U1118 ( .A(n9), .B(n1353), .C(n6), .D(n1352), .Z(n1066) );
  COND2X1 U1119 ( .A(n9), .B(n1354), .C(n6), .D(n1353), .Z(n1067) );
  COND2X1 U1120 ( .A(n9), .B(n1355), .C(n6), .D(n1354), .Z(n1068) );
  COND2X1 U1122 ( .A(n9), .B(n1357), .C(n6), .D(n1356), .Z(n1070) );
  COND2X1 U1123 ( .A(n9), .B(n1358), .C(n6), .D(n1357), .Z(n1071) );
  COND2X1 U1124 ( .A(n9), .B(n1359), .C(n6), .D(n1358), .Z(n1072) );
  COND2X1 U1125 ( .A(n9), .B(n1360), .C(n6), .D(n1359), .Z(n1073) );
  COND2X1 U1126 ( .A(n9), .B(n1361), .C(n6), .D(n1360), .Z(n1074) );
  COND2X1 U1127 ( .A(n9), .B(n1362), .C(n6), .D(n1361), .Z(n1075) );
  COND2X1 U1128 ( .A(n9), .B(n1363), .C(n6), .D(n1362), .Z(n1076) );
  COND2X1 U1129 ( .A(n9), .B(n1364), .C(n6), .D(n1363), .Z(n1077) );
  COND2X1 U1130 ( .A(n9), .B(n1365), .C(n6), .D(n1364), .Z(n1078) );
  COND2X1 U1131 ( .A(n9), .B(n1366), .C(n6), .D(n1365), .Z(n1079) );
  COND2X1 U1132 ( .A(n9), .B(n1367), .C(n6), .D(n1366), .Z(n1080) );
  COND2X1 U1133 ( .A(n9), .B(n1368), .C(n6), .D(n1367), .Z(n1081) );
  COND2X1 U1135 ( .A(n9), .B(n1370), .C(n6), .D(n1369), .Z(n1083) );
  COND2X1 U1136 ( .A(n9), .B(n1371), .C(n6), .D(n1370), .Z(n1084) );
  COND2X1 U1137 ( .A(n9), .B(n1372), .C(n6), .D(n1371), .Z(n1085) );
  CEOX2 U1260 ( .A(a[2]), .B(n2229), .Z(n1420) );
  CEOX2 U1263 ( .A(a[0]), .B(n2221), .Z(n1421) );
  CFD1QXL clk_r_REG14_S1 ( .D(n254), .CP(n2183), .Q(n2181) );
  CFD1QXL clk_r_REG4_S1 ( .D(n279), .CP(n2183), .Q(n2161) );
  CFD1QXL clk_r_REG6_S1 ( .D(n138), .CP(n2183), .Q(n2174) );
  CFD1QXL clk_r_REG1_S1 ( .D(n295), .CP(n2183), .Q(n2167) );
  CFD1QXL clk_r_REG163_S1 ( .D(n845), .CP(n2183), .Q(n2038) );
  CFD1QXL clk_r_REG123_S1 ( .D(n947), .CP(n2183), .Q(n2051) );
  CFD1QXL clk_r_REG102_S1 ( .D(n397), .CP(n2183), .Q(n2159) );
  CFD1QXL clk_r_REG132_S1 ( .D(n925), .CP(n2183), .Q(n2041) );
  CFD1QXL clk_r_REG150_S1 ( .D(n887), .CP(n2183), .Q(n2036) );
  CFD1QXL clk_r_REG144_S1 ( .D(n905), .CP(n2183), .Q(n2058) );
  CFD1QXL clk_r_REG101_S1 ( .D(n1055), .CP(n2183), .Q(n2047) );
  CFD1QXL clk_r_REG103_S1 ( .D(n398), .CP(n2183), .Q(n2158) );
  CFD1QXL clk_r_REG33_S1 ( .D(n641), .CP(n2183), .Q(n2102) );
  CFD1QXL clk_r_REG21_S1 ( .D(n659), .CP(n2183), .Q(n2095) );
  CFD1QXL clk_r_REG71_S1 ( .D(n609), .CP(n2183), .Q(n2116) );
  CFD1QXL clk_r_REG117_S1 ( .D(n454), .CP(n2183), .Q(n2150) );
  CFD1QXL clk_r_REG60_S1 ( .D(n596), .CP(n2183), .Q(n2119) );
  CFD1QXL clk_r_REG126_S1 ( .D(n526), .CP(n2183), .Q(n2139) );
  CFD1QXL clk_r_REG137_S1 ( .D(n612), .CP(n2183), .Q(n2169) );
  CFD1QXL clk_r_REG120_S1 ( .D(n550), .CP(n2183), .Q(n2135) );
  CFD1QXL clk_r_REG49_S1 ( .D(n508), .CP(n2183), .Q(n2143) );
  CFD1QXL clk_r_REG54_S1 ( .D(n625), .CP(n2183), .Q(n2110) );
  CFD1QXL clk_r_REG135_S1 ( .D(n926), .CP(n2183), .Q(n2042) );
  CFD1QXL clk_r_REG109_S1 ( .D(n373), .CP(n2183), .Q(n2166) );
  CFD1QXL clk_r_REG159_S1 ( .D(n857), .CP(n2183), .Q(n2064) );
  CFD1QXL clk_r_REG167_S1 ( .D(n799), .CP(n2183), .Q(n2088) );
  CFD1QXL clk_r_REG142_S1 ( .D(n815), .CP(n2183), .Q(n2087) );
  CFD1QXL clk_r_REG99_S1 ( .D(n817), .CP(n2183), .Q(n2086) );
  CFD1QXL clk_r_REG9_S1 ( .D(n272), .CP(n2183), .Q(n2177) );
  CFD1QXL clk_r_REG30_S1 ( .D(n423), .CP(n2183), .Q(n2153) );
  CFD1QXL clk_r_REG47_S1 ( .D(n522), .CP(n2183), .Q(n2141) );
  CFD1QXL clk_r_REG18_S1 ( .D(n657), .CP(n2183), .Q(n2097) );
  CFD1QXL clk_r_REG20_S1 ( .D(n673), .CP(n2183), .Q(n2090) );
  CFD1QXL clk_r_REG113_S1 ( .D(n478), .CP(n2183), .Q(n2148) );
  CFD1QXL clk_r_REG134_S1 ( .D(n592), .CP(n2183), .Q(n2123) );
  CFD1QXL clk_r_REG81_S1 ( .D(n501), .CP(n2183), .Q(net171643) );
  CFD1QXL clk_r_REG115_S1 ( .D(n504), .CP(n2183), .Q(n2145) );
  CFD1QXL clk_r_REG112_S1 ( .D(n477), .CP(n2183), .Q(n2149) );
  CFD1QXL clk_r_REG24_S1 ( .D(n614), .CP(n2183), .Q(n2113) );
  CFD1QXL clk_r_REG29_S1 ( .D(n1611), .CP(n2183), .Q(n2165) );
  CFD1QXL clk_r_REG130_S1 ( .D(n427), .CP(n2183), .Q(net171635) );
  CFD1QXL clk_r_REG45_S1 ( .D(n531), .CP(n2183), .Q(n2138) );
  CFD1QXL clk_r_REG67_S1 ( .D(n486), .CP(n2183), .Q(n2164) );
  CFD1QXL clk_r_REG35_S1 ( .D(n645), .CP(n2183), .Q(n2100) );
  CFD1QXL clk_r_REG46_S1 ( .D(n521), .CP(n2183), .Q(n2142) );
  CFD1QXL clk_r_REG73_S1 ( .D(n576), .CP(n2183), .Q(n2125) );
  CFD1QXL clk_r_REG52_S1 ( .D(n628), .CP(n2183), .Q(n2107) );
  CFD1QXL clk_r_REG36_S1 ( .D(n646), .CP(n2183), .Q(n2099) );
  CFD1QXL clk_r_REG39_S1 ( .D(n569), .CP(n2183), .Q(n2129) );
  CFD1QXL clk_r_REG41_S1 ( .D(n547), .CP(n2183), .Q(n2137) );
  CFD1QXL clk_r_REG66_S1 ( .D(n485), .CP(n2183), .Q(net171503) );
  CFD1QXL clk_r_REG111_S1 ( .D(n452), .CP(n2183), .Q(n2151) );
  CFD1QXL clk_r_REG118_S1 ( .D(n998), .CP(n2183), .Q(n2034) );
  CFD1QXL clk_r_REG125_S1 ( .D(n525), .CP(n2183), .Q(n2140) );
  CFD1QXL clk_r_REG65_S1 ( .D(n630), .CP(n2183), .Q(n2105) );
  CFD1QXL clk_r_REG51_S1 ( .D(n627), .CP(n2183), .Q(n2108) );
  CFD1QXL clk_r_REG133_S1 ( .D(n591), .CP(n2183), .Q(n2124) );
  CFD1QXL clk_r_REG121_S1 ( .D(n571), .CP(n2183), .Q(n2127) );
  CFD1QXL clk_r_REG8_S1 ( .D(n276), .CP(n2183), .Q(n2176) );
  CFD1QXL clk_r_REG16_S1 ( .D(n671), .CP(n2183), .Q(n2092) );
  CFD1QXL clk_r_REG15_S1 ( .D(n687), .CP(n2183), .Q(n2089) );
  CFD1QXL clk_r_REG10_S1 ( .D(n271), .CP(n2183), .Q(n2178) );
  CFD1QXL clk_r_REG7_S1 ( .D(n277), .CP(n2183), .Q(n2175) );
  CFD1QX2 clk_r_REG162_S1 ( .D(n913), .CP(n2183), .Q(n2052) );
  CFD1QX2 clk_r_REG153_S1 ( .D(n955), .CP(n2183), .Q(n2049) );
  CFD1QX2 clk_r_REG171_S1 ( .D(n800), .CP(n2183), .Q(net171759) );
  CFD1QX2 clk_r_REG58_S1 ( .D(n848), .CP(n2183), .Q(n2066) );
  CFD1QX2 clk_r_REG164_S1 ( .D(n826), .CP(n2183), .Q(n2170) );
  CFD1QX2 clk_r_REG43_S1 ( .D(n860), .CP(n2183), .Q(n2063) );
  CFD1QX2 clk_r_REG139_S1 ( .D(n833), .CP(n2183), .Q(n2071) );
  CFD1QX2 clk_r_REG122_S1 ( .D(n572), .CP(n2183), .Q(n2126) );
  CFD1QX2 clk_r_REG106_S1 ( .D(n824), .CP(n2183), .Q(n2080) );
  CFD1QX2 clk_r_REG161_S1 ( .D(n874), .CP(n2183), .Q(n2060) );
  CFD1QX2 clk_r_REG170_S1 ( .D(n801), .CP(n2183), .Q(net171708) );
  CFD1QX2 clk_r_REG44_S1 ( .D(n861), .CP(n2183), .Q(n2062) );
  CFD1QX2 clk_r_REG55_S1 ( .D(n626), .CP(n2183), .Q(n2109) );
  CFD1QX2 clk_r_REG37_S1 ( .D(n553), .CP(n2183), .Q(n2133) );
  CFD1QX2 clk_r_REG97_S1 ( .D(n831), .CP(n2183), .Q(n2073) );
  CFD1QX2 clk_r_REG119_S1 ( .D(n1061), .CP(n2183), .Q(n2045) );
  CFD1QX1 clk_r_REG78_S1 ( .D(n555), .CP(n2183), .Q(n2131) );
  CFD1QX2 clk_r_REG143_S1 ( .D(n951), .CP(n2183), .Q(n2040) );
  CFD1QX2 clk_r_REG140_S1 ( .D(n825), .CP(n2183), .Q(n2079) );
  CFD1QX2 clk_r_REG76_S1 ( .D(n828), .CP(n2183), .Q(n2076) );
  CFD1QX1 clk_r_REG80_S1 ( .D(n534), .CP(n2183), .Q(n2163) );
  CFD1QX2 clk_r_REG84_S1 ( .D(n829), .CP(n2183), .Q(n2075) );
  CFD1QX1 clk_r_REG12_S1 ( .D(n2013), .CP(n2183), .Q(n2182) );
  CFD1QX1 clk_r_REG70_S1 ( .D(n617), .CP(n2183), .Q(n2162) );
  CFD1QX2 clk_r_REG69_S1 ( .D(n827), .CP(n2183), .Q(n2077) );
  CFD1QX2 clk_r_REG88_S1 ( .D(n615), .CP(n2183), .Q(n2112) );
  CFD1QX2 clk_r_REG11_S1 ( .D(n267), .CP(n2183), .Q(n2179) );
  CFD1QX2 clk_r_REG31_S1 ( .D(n424), .CP(n2183), .Q(net171634) );
  CFD1QX2 clk_r_REG13_S1 ( .D(n255), .CP(n2183), .Q(n2180) );
  CFD1QX1 clk_r_REG42_S1 ( .D(n548), .CP(n2183), .Q(n2136) );
  CFD1QX1 clk_r_REG87_S1 ( .D(n652), .CP(n2183), .Q(n2098) );
  CFD1QX1 clk_r_REG50_S1 ( .D(n650), .CP(n2183), .Q(n2039) );
  CFD1QX1 clk_r_REG23_S1 ( .D(n613), .CP(n2183), .Q(n2114) );
  CFD1QX4 clk_r_REG68_S1 ( .D(n837), .CP(n2183), .Q(net171723) );
  CFD1QX2 clk_r_REG57_S1 ( .D(n633), .CP(n2183), .Q(n2103) );
  CFD1QX2 clk_r_REG94_S1 ( .D(n597), .CP(n2183), .Q(n2118) );
  CFD1QX1 clk_r_REG53_S1 ( .D(n631), .CP(n2183), .Q(n2104) );
  CFD1QX2 clk_r_REG89_S1 ( .D(n616), .CP(n2183), .Q(n2111) );
  CFD1QX2 clk_r_REG59_S1 ( .D(n595), .CP(n2183), .Q(n2120) );
  CFD1QX2 clk_r_REG98_S1 ( .D(n823), .CP(n2183), .Q(n2081) );
  CFD1QX1 clk_r_REG146_S1 ( .D(n906), .CP(n2183), .Q(n2057) );
  CFD1QX4 clk_r_REG91_S1 ( .D(n840), .CP(n2183), .Q(n2068) );
  CFD1QX1 clk_r_REG61_S1 ( .D(n552), .CP(n2183), .Q(n2134) );
  CFD1QX4 clk_r_REG157_S1 ( .D(n911), .CP(n2183), .Q(n2053) );
  CFD1QX2 clk_r_REG148_S1 ( .D(n953), .CP(n2183), .Q(n2050) );
  CFD1QX1 clk_r_REG108_S1 ( .D(n1057), .CP(n2183), .Q(n2046) );
  CFD1QX1 clk_r_REG124_S1 ( .D(n973), .CP(n2183), .Q(n2048) );
  CFD1QX2 clk_r_REG96_S1 ( .D(n841), .CP(n2183), .Q(n2067) );
  CFD1QX1 clk_r_REG38_S1 ( .D(n554), .CP(n2183), .Q(n2132) );
  CFD1QX2 clk_r_REG105_S1 ( .D(n832), .CP(n2183), .Q(n2072) );
  CFD1QX2 clk_r_REG158_S1 ( .D(n891), .CP(n2183), .Q(n2037) );
  CFD1QX4 clk_r_REG74_S1 ( .D(n850), .CP(n2183), .Q(n2065) );
  CFD1QX4 clk_r_REG155_S1 ( .D(n910), .CP(n2183), .Q(n2054) );
  CFD1QX1 clk_r_REG145_S1 ( .D(n927), .CP(n2183), .Q(n2043) );
  CFD1QX4 clk_r_REG169_S1 ( .D(n802), .CP(n2183), .Q(n2078) );
  CFD1QX1 clk_r_REG131_S1 ( .D(n428), .CP(n2183), .Q(n2152) );
  CFD1QX4 clk_r_REG151_S1 ( .D(n929), .CP(n2183), .Q(net171752) );
  CFD1QX2 clk_r_REG165_S1 ( .D(n820), .CP(n2183), .Q(n2171) );
  CFD1QX2 clk_r_REG48_S1 ( .D(n507), .CP(n2183), .Q(n2144) );
  CFD1QX2 clk_r_REG92_S1 ( .D(n830), .CP(n2183), .Q(n2074) );
  CFD1QX1 clk_r_REG64_S1 ( .D(n629), .CP(n2183), .Q(n2106) );
  CFA1X1 U428 ( .A(n470), .B(n491), .CI(n468), .CO(n463), .S(n464) );
  CFA1X1 U427 ( .A(n466), .B(n464), .CI(n489), .CO(n461), .S(n462) );
  CFA1X1 U388 ( .A(n390), .B(n413), .CI(n415), .CO(n383), .S(n384) );
  CFA1X1 U403 ( .A(n445), .B(n422), .CI(n420), .CO(n413), .S(n414) );
  CFA1X1 U386 ( .A(n384), .B(n382), .CI(n409), .CO(n379), .S(n380) );
  CFA1X1 U401 ( .A(n416), .B(n439), .CI(n414), .CO(n409), .S(n410) );
  CFA1X1 U400 ( .A(net179910), .B(n410), .CI(n437), .CO(n407), .S(n408) );
  CFD1QX1 clk_r_REG114_S1 ( .D(n503), .CP(n2183), .Q(n2146) );
  CFD1QX4 clk_r_REG152_S1 ( .D(n908), .CP(n2183), .Q(n2056) );
  CFD1QXL clk_r_REG5_S1 ( .D(n140), .CP(n2183), .Q(n2173) );
  CFD1QXL clk_r_REG22_S1 ( .D(n660), .CP(n2183), .Q(n2094) );
  CFD1QXL clk_r_REG128_S1 ( .D(n399), .CP(n2183), .Q(n2157) );
  CFD1QX2 clk_r_REG107_S1 ( .D(n818), .CP(n2183), .Q(n2085) );
  CFD1QX2 clk_r_REG19_S1 ( .D(n658), .CP(n2183), .Q(n2096) );
  CFD1QX2 clk_r_REG85_S1 ( .D(n821), .CP(n2183), .Q(n2083) );
  CFD1QX2 clk_r_REG27_S1 ( .D(n405), .CP(n2183), .Q(n2155) );
  CFD1QX1 clk_r_REG34_S1 ( .D(n642), .CP(n2183), .Q(n2101) );
  CFD1QX1 clk_r_REG25_S1 ( .D(n593), .CP(n2183), .Q(n2122) );
  CFD1QX2 clk_r_REG72_S1 ( .D(n610), .CP(n2183), .Q(n2115) );
  CFD1QX2 clk_r_REG138_S1 ( .D(n611), .CP(n2183), .Q(n2160) );
  CFD1QX2 clk_r_REG40_S1 ( .D(n570), .CP(n2183), .Q(n2128) );
  CFD1QX2 clk_r_REG154_S1 ( .D(n909), .CP(n2183), .Q(n2055) );
  CFD1QX2 clk_r_REG156_S1 ( .D(n872), .CP(n2183), .Q(n2061) );
  CFD1QX4 clk_r_REG160_S1 ( .D(n892), .CP(n2183), .Q(n2059) );
  CFD1QX1 clk_r_REG79_S1 ( .D(n556), .CP(n2183), .Q(n2130) );
  CFD1QX2 clk_r_REG93_S1 ( .D(n822), .CP(n2183), .Q(n2082) );
  CFD1QX2 clk_r_REG129_S1 ( .D(n400), .CP(n2183), .Q(n2156) );
  CFD1QX1 clk_r_REG82_S1 ( .D(n502), .CP(n2183), .Q(n2147) );
  CFD1QX2 clk_r_REG168_S1 ( .D(n803), .CP(n2183), .Q(n2070) );
  CFD1QXL clk_r_REG17_S1 ( .D(n672), .CP(n2183), .Q(n2091) );
  CFD1QX2 clk_r_REG83_S1 ( .D(n839), .CP(n2183), .Q(net171725) );
  CFD1QX2 clk_r_REG62_S1 ( .D(n665), .CP(n2183), .Q(n2093) );
  CFD1QX1 clk_r_REG127_S1 ( .D(n1001), .CP(n2183), .Q(n2035) );
  CFD1QX2 clk_r_REG28_S1 ( .D(n406), .CP(n2183), .Q(n2154) );
  CFD1QX4 clk_r_REG147_S1 ( .D(n928), .CP(n2183), .Q(n2044) );
  CFD1QX4 clk_r_REG75_S1 ( .D(n838), .CP(n2183), .Q(n2069) );
  CFD1QX4 clk_r_REG149_S1 ( .D(n907), .CP(n2183), .Q(net171738) );
  CFD1QX2 clk_r_REG95_S1 ( .D(n598), .CP(n2183), .Q(n2117) );
  CFD1QX1 clk_r_REG26_S1 ( .D(n594), .CP(n2183), .Q(n2121) );
  CFD1QX2 clk_r_REG2_S1 ( .D(n284), .CP(n2183), .Q(n2168) );
  CFD1QX2 clk_r_REG141_S1 ( .D(n819), .CP(n2183), .Q(n2084) );
  CFD1QX2 clk_r_REG32_S1 ( .D(n378), .CP(n2183), .Q(n2172) );
  CFD1QX2 clk_r_REG116_S1 ( .D(n453), .CP(n2183), .Q(net171639) );
  CFD1QX4 clk_r_REG110_S1 ( .D(n451), .CP(n2183), .Q(net171637) );
  CND2X2 U1267 ( .A(n458), .B(n2150), .Z(n1654) );
  CENX2 U1268 ( .A(net171637), .B(net171639), .Z(net182724) );
  CIVX1 U1269 ( .A(n229), .Z(n227) );
  CND2X2 U1270 ( .A(n2059), .B(n2054), .Z(n1920) );
  CNR2X1 U1271 ( .A(net179493), .B(n435), .Z(n1690) );
  CEOXL U1272 ( .A(n1953), .B(n500), .Z(n494) );
  CND2X2 U1273 ( .A(n500), .B(n2142), .Z(n1955) );
  CND2X2 U1274 ( .A(n2060), .B(n2044), .Z(n1721) );
  CEO3X1 U1275 ( .A(n2074), .B(n2044), .C(n2060), .Z(n458) );
  CENX1 U1276 ( .A(net33482), .B(n2002), .Z(n1182) );
  CENXL U1277 ( .A(n2221), .B(n1388), .Z(n1355) );
  CENXL U1278 ( .A(n2221), .B(n1389), .Z(n1356) );
  CENXL U1279 ( .A(n2221), .B(n2209), .Z(n1360) );
  CENXL U1280 ( .A(net33080), .B(n2221), .Z(n1372) );
  CENXL U1281 ( .A(n2221), .B(n2210), .Z(n1359) );
  CENXL U1282 ( .A(n2221), .B(n2212), .Z(n1357) );
  CENXL U1283 ( .A(n2221), .B(n2211), .Z(n1358) );
  CNIVX3 U1284 ( .A(n63), .Z(n2002) );
  CND2X1 U1285 ( .A(n1411), .B(n89), .Z(n91) );
  CND2X4 U1286 ( .A(n1772), .B(n1773), .Z(n1411) );
  CIVX2 U1287 ( .A(n1780), .Z(n1765) );
  CEO3X1 U1288 ( .A(net171634), .B(n449), .C(n447), .Z(n1779) );
  CNIVX4 U1289 ( .A(n93), .Z(n1963) );
  CND2X4 U1290 ( .A(n1411), .B(n89), .Z(n1964) );
  CND2X1 U1291 ( .A(n2171), .B(n2069), .Z(n1930) );
  CND2X1 U1292 ( .A(n2171), .B(n2066), .Z(n1931) );
  CEOX1 U1293 ( .A(n1737), .B(n2062), .Z(n482) );
  CEOX2 U1294 ( .A(n2055), .B(n2073), .Z(n1737) );
  CND2X2 U1295 ( .A(n2072), .B(n2054), .Z(n1919) );
  CNR2X1 U1296 ( .A(net179834), .B(n487), .Z(n1937) );
  CENX1 U1297 ( .A(n2201), .B(n1755), .Z(n1692) );
  COR2XL U1298 ( .A(n2001), .B(n2000), .Z(n1543) );
  CENX2 U1299 ( .A(n873), .B(n1544), .Z(n434) );
  CNR2X2 U1300 ( .A(n2001), .B(n2000), .Z(n1544) );
  CEO3X1 U1301 ( .A(n2074), .B(n2044), .C(n2060), .Z(n1545) );
  CND2X1 U1302 ( .A(n2074), .B(n2060), .Z(n1719) );
  CND2X1 U1303 ( .A(n2074), .B(n2044), .Z(n1720) );
  CEOX2 U1304 ( .A(n450), .B(n471), .Z(n1546) );
  CEOX2 U1305 ( .A(n448), .B(n1546), .Z(n442) );
  CND2X1 U1306 ( .A(n448), .B(n471), .Z(n1547) );
  CND2X1 U1307 ( .A(n448), .B(n450), .Z(n1548) );
  CND2X1 U1308 ( .A(n471), .B(n450), .Z(n1549) );
  CND3X2 U1309 ( .A(n1547), .B(n1548), .C(n1549), .Z(n441) );
  CENX1 U1310 ( .A(n1556), .B(n430), .Z(n1741) );
  CND2XL U1311 ( .A(n430), .B(n2152), .Z(n1744) );
  CND2XL U1312 ( .A(n426), .B(n430), .Z(n1742) );
  CND2XL U1313 ( .A(n426), .B(n2152), .Z(n1743) );
  CND2X1 U1314 ( .A(n493), .B(n495), .Z(n1604) );
  CHA1X1 U1315 ( .A(n895), .B(n865), .CO(n577), .S(n578) );
  CIVXL U1316 ( .A(n463), .Z(n1550) );
  CIVXL U1317 ( .A(n1550), .Z(n1551) );
  CIVX4 U1318 ( .A(n2033), .Z(n2184) );
  CENXL U1319 ( .A(n1552), .B(n843), .Z(n572) );
  CENX1 U1320 ( .A(n1063), .B(n979), .Z(n1552) );
  CENX1 U1321 ( .A(n689), .B(n676), .Z(n1615) );
  CENX1 U1322 ( .A(n1553), .B(n992), .Z(n766) );
  CENX1 U1323 ( .A(n946), .B(n968), .Z(n1553) );
  CND2XL U1324 ( .A(n647), .B(n651), .Z(n1651) );
  CEOXL U1325 ( .A(n1648), .B(n651), .Z(n628) );
  CND2XL U1326 ( .A(n551), .B(n549), .Z(n1888) );
  CEOXL U1327 ( .A(n549), .B(n551), .Z(n1885) );
  CIVXL U1328 ( .A(n89), .Z(n1554) );
  CIVXL U1329 ( .A(n1554), .Z(n1555) );
  CIVX20 U1330 ( .A(n2152), .Z(n1556) );
  CIVX2 U1331 ( .A(n1804), .Z(n1805) );
  COND2X1 U1332 ( .A(n107), .B(n1098), .C(n105), .D(n1097), .Z(n824) );
  CHA1X1 U1333 ( .A(n897), .B(n867), .CO(n617), .S(n618) );
  CND2X1 U1334 ( .A(net178620), .B(n156), .Z(n120) );
  COND2XL U1335 ( .A(n1095), .B(n107), .C(n105), .D(n1094), .Z(n821) );
  CND2XL U1336 ( .A(n1777), .B(n1776), .Z(n1558) );
  CND2X2 U1337 ( .A(n1777), .B(n1776), .Z(n114) );
  CNIVX4 U1338 ( .A(n66), .Z(n1607) );
  CENX2 U1339 ( .A(n1944), .B(n1557), .Z(n676) );
  CEN3X2 U1340 ( .A(n919), .B(n985), .C(n1613), .Z(n1557) );
  CFA1XL U1341 ( .A(n844), .B(n854), .CI(n866), .CO(n597), .S(n598) );
  CND3X1 U1342 ( .A(n1645), .B(n1646), .C(n1647), .Z(n651) );
  CIVX2 U1343 ( .A(n109), .Z(n1774) );
  CIVX3 U1344 ( .A(n109), .Z(n1432) );
  CNR2IX2 U1345 ( .B(net33082), .A(n114), .Z(n816) );
  CANR1X1 U1346 ( .A(n185), .B(n1662), .C(n173), .Z(n171) );
  CENXL U1347 ( .A(net33482), .B(n113), .Z(n1086) );
  CEOXL U1348 ( .A(a[30]), .B(a[31]), .Z(n1406) );
  CND2XL U1349 ( .A(n114), .B(n1406), .Z(n115) );
  CIVX2 U1350 ( .A(n2230), .Z(n2227) );
  CIVX2 U1351 ( .A(n2230), .Z(n2226) );
  CIVX3 U1352 ( .A(n2230), .Z(n2225) );
  CIVX3 U1353 ( .A(n2230), .Z(n2228) );
  CIVX3 U1354 ( .A(n2230), .Z(n2224) );
  CIVX8 U1355 ( .A(n12), .Z(n2230) );
  CIVX2 U1356 ( .A(n2002), .Z(n1559) );
  CIVX3 U1357 ( .A(n1559), .Z(n1560) );
  CNIVX4 U1358 ( .A(n1397), .Z(n2206) );
  CNIVX1 U1359 ( .A(n1745), .Z(n1561) );
  CENXL U1360 ( .A(n1562), .B(n816), .Z(n406) );
  CENX1 U1361 ( .A(n846), .B(n836), .Z(n1562) );
  CND2X1 U1362 ( .A(n436), .B(n461), .Z(net179954) );
  CNR2X2 U1363 ( .A(net179805), .B(n461), .Z(n167) );
  CND2XL U1364 ( .A(n2149), .B(n1699), .Z(n1935) );
  CND3X1 U1365 ( .A(n1933), .B(n1934), .C(n1935), .Z(n447) );
  CIVX1 U1366 ( .A(n156), .Z(n154) );
  CEOX1 U1367 ( .A(n723), .B(n712), .Z(n1563) );
  CEOX1 U1368 ( .A(n1563), .B(n721), .Z(n706) );
  CND2XL U1369 ( .A(n721), .B(n712), .Z(n1564) );
  CND2XL U1370 ( .A(n721), .B(n723), .Z(n1565) );
  CND2XL U1371 ( .A(n712), .B(n723), .Z(n1566) );
  CND3X1 U1372 ( .A(n1564), .B(n1565), .C(n1566), .Z(n705) );
  CFA1XL U1373 ( .A(n964), .B(n1072), .CI(n1042), .CO(n723), .S(n724) );
  CENXL U1374 ( .A(net33482), .B(n109), .Z(n1091) );
  CND2IXL U1375 ( .B(n1963), .A(n1993), .Z(n1989) );
  CEO3X2 U1376 ( .A(n2171), .B(n2069), .C(n2066), .Z(n460) );
  CND2XL U1377 ( .A(n649), .B(n651), .Z(n1650) );
  CND2XL U1378 ( .A(n899), .B(n805), .Z(n1646) );
  CND2XL U1379 ( .A(n869), .B(n805), .Z(n1647) );
  CND2XL U1380 ( .A(n479), .B(n1699), .Z(n1934) );
  CND2XL U1381 ( .A(n479), .B(n2149), .Z(n1933) );
  CEO3X2 U1382 ( .A(n748), .B(n753), .C(n746), .Z(n742) );
  CEOX2 U1383 ( .A(n751), .B(n744), .Z(n1567) );
  CEOX2 U1384 ( .A(n1567), .B(n742), .Z(n740) );
  CND2XL U1385 ( .A(n748), .B(n753), .Z(n1568) );
  CND2XL U1386 ( .A(n748), .B(n746), .Z(n1569) );
  CND2XL U1387 ( .A(n753), .B(n746), .Z(n1570) );
  CND3X1 U1388 ( .A(n1568), .B(n1569), .C(n1570), .Z(n741) );
  CND2XL U1389 ( .A(n751), .B(n744), .Z(n1571) );
  CND2XL U1390 ( .A(n751), .B(n742), .Z(n1572) );
  CND2XL U1391 ( .A(n744), .B(n742), .Z(n1573) );
  CND3XL U1392 ( .A(n1571), .B(n1572), .C(n1573), .Z(n739) );
  CEOX1 U1393 ( .A(n1017), .B(n991), .Z(n1574) );
  CEOX2 U1394 ( .A(n1574), .B(n758), .Z(n754) );
  CND2XL U1395 ( .A(n758), .B(n991), .Z(n1575) );
  CND2XL U1396 ( .A(n758), .B(n1017), .Z(n1576) );
  CND2XL U1397 ( .A(n991), .B(n1017), .Z(n1577) );
  CND3X1 U1398 ( .A(n1575), .B(n1576), .C(n1577), .Z(n753) );
  CIVXL U1399 ( .A(n1545), .Z(n1578) );
  CIVXL U1400 ( .A(n1578), .Z(n1579) );
  CIVX4 U1401 ( .A(n55), .Z(n2256) );
  CIVXL U1402 ( .A(n459), .Z(n1580) );
  CIVXL U1403 ( .A(n1580), .Z(n1581) );
  CEO3X2 U1404 ( .A(n420), .B(net184228), .C(n1657), .Z(net179947) );
  CND2X1 U1405 ( .A(a[28]), .B(n1774), .Z(n1584) );
  CND2X2 U1406 ( .A(n1582), .B(n1583), .Z(n1585) );
  CND2X2 U1407 ( .A(n1584), .B(n1585), .Z(n1407) );
  CIVXL U1408 ( .A(a[28]), .Z(n1582) );
  CIVX2 U1409 ( .A(n1774), .Z(n1583) );
  CEO3X2 U1410 ( .A(n517), .B(n515), .C(n494), .Z(n490) );
  CEOX2 U1411 ( .A(n492), .B(n513), .Z(n1586) );
  CEOX1 U1412 ( .A(n1586), .B(n490), .Z(n488) );
  CND2XL U1413 ( .A(n517), .B(n515), .Z(n1587) );
  CND2XL U1414 ( .A(n517), .B(n494), .Z(n1588) );
  CND2XL U1415 ( .A(n515), .B(n494), .Z(n1589) );
  CND3X1 U1416 ( .A(n1587), .B(n1588), .C(n1589), .Z(n489) );
  CND2XL U1417 ( .A(n492), .B(n513), .Z(n1590) );
  CND2X1 U1418 ( .A(n492), .B(n490), .Z(n1591) );
  CND2X1 U1419 ( .A(n513), .B(n490), .Z(n1592) );
  CND3X2 U1420 ( .A(n1590), .B(n1591), .C(n1592), .Z(n487) );
  CEOX1 U1421 ( .A(n2141), .B(n543), .Z(n1593) );
  CEOX2 U1422 ( .A(n1593), .B(n520), .Z(n516) );
  CND2X1 U1423 ( .A(n520), .B(n543), .Z(n1594) );
  CND2X1 U1424 ( .A(n520), .B(n2141), .Z(n1595) );
  CND2X1 U1425 ( .A(n543), .B(n2141), .Z(n1596) );
  CND3X2 U1426 ( .A(n1594), .B(n1595), .C(n1596), .Z(n515) );
  CENX1 U1427 ( .A(n528), .B(n1823), .Z(n520) );
  CIVXL U1428 ( .A(n445), .Z(n1656) );
  CNR2XL U1429 ( .A(n488), .B(n511), .Z(n1597) );
  CND2X1 U1430 ( .A(n2053), .B(n2078), .Z(n1600) );
  CND2X2 U1431 ( .A(n1598), .B(n1599), .Z(n1601) );
  CND2X2 U1432 ( .A(n1600), .B(n1601), .Z(n1756) );
  CIVX2 U1433 ( .A(n2053), .Z(n1598) );
  CIVX3 U1434 ( .A(n2078), .Z(n1599) );
  CEOX2 U1435 ( .A(n495), .B(n472), .Z(n1602) );
  CEOX2 U1436 ( .A(n1602), .B(n493), .Z(n466) );
  CND2XL U1437 ( .A(n493), .B(n472), .Z(n1603) );
  CND2XL U1438 ( .A(n472), .B(n495), .Z(n1605) );
  CND3X2 U1439 ( .A(n1603), .B(n1604), .C(n1605), .Z(n465) );
  CEO3X2 U1440 ( .A(n1793), .B(n480), .C(n1798), .Z(n472) );
  CEO3X1 U1441 ( .A(n444), .B(n442), .C(n465), .Z(net179996) );
  CND3X1 U1442 ( .A(n1716), .B(n1717), .C(n1718), .Z(n495) );
  CENX2 U1443 ( .A(n1851), .B(n460), .Z(n448) );
  CND2X1 U1444 ( .A(n2035), .B(n2164), .Z(n1838) );
  CEO3X1 U1445 ( .A(n2035), .B(n509), .C(n2164), .Z(n476) );
  CNR2X1 U1446 ( .A(n1123), .B(n89), .Z(n2001) );
  COND2X1 U1447 ( .A(n1964), .B(n1132), .C(n89), .D(n1131), .Z(n855) );
  CENX1 U1448 ( .A(n2068), .B(n2065), .Z(n1992) );
  CIVX4 U1449 ( .A(n21), .Z(n2237) );
  CNR2IX1 U1450 ( .B(n1684), .A(n1677), .Z(n1681) );
  CANR1XL U1451 ( .A(n425), .B(n1677), .C(net171635), .Z(n1682) );
  CEOX1 U1452 ( .A(n1913), .B(n699), .Z(n678) );
  CND2X1 U1453 ( .A(n2068), .B(n1701), .Z(n1702) );
  CND2X1 U1454 ( .A(n1700), .B(n2065), .Z(n1703) );
  CENX1 U1455 ( .A(n2247), .B(net33480), .Z(n1250) );
  CND2X1 U1456 ( .A(n2037), .B(n2040), .Z(n1749) );
  CND2X1 U1457 ( .A(n2037), .B(n2079), .Z(n1750) );
  CND2X1 U1458 ( .A(n2040), .B(n2079), .Z(n1751) );
  CFA1X1 U1459 ( .A(n1018), .B(n1076), .CI(n1046), .CO(n763), .S(n764) );
  CND2X1 U1460 ( .A(net171723), .B(n1687), .Z(n1680) );
  CNR2X1 U1461 ( .A(net171723), .B(n1687), .Z(n1679) );
  CND2X1 U1462 ( .A(n1728), .B(n1729), .Z(n1761) );
  CND2X1 U1463 ( .A(n1726), .B(n1727), .Z(n1729) );
  CND2X1 U1464 ( .A(n607), .B(n605), .Z(n1845) );
  CND2X1 U1465 ( .A(n605), .B(n590), .Z(n1847) );
  CND3X1 U1466 ( .A(n1837), .B(n1838), .C(n1839), .Z(n475) );
  CND3X1 U1467 ( .A(n1896), .B(n1897), .C(n1898), .Z(n519) );
  CEOX1 U1468 ( .A(n1670), .B(n510), .Z(n498) );
  CENX1 U1469 ( .A(n1867), .B(n545), .Z(n518) );
  CIVX2 U1470 ( .A(n39), .Z(n2250) );
  COND2XL U1471 ( .A(n1148), .B(n1864), .C(n1978), .D(n84), .Z(n805) );
  CND3X1 U1472 ( .A(n1852), .B(n1853), .C(n1854), .Z(n683) );
  CIVX4 U1473 ( .A(n2029), .Z(n33) );
  CNIVX4 U1474 ( .A(n116), .Z(net33082) );
  CNR2IX1 U1475 ( .B(net33082), .A(n95), .Z(n844) );
  CND2X1 U1476 ( .A(n1976), .B(n1977), .Z(n804) );
  CAN2X1 U1477 ( .A(n1802), .B(n151), .Z(net179380) );
  CIVXL U1478 ( .A(n39), .Z(n2251) );
  CIVX1 U1479 ( .A(n2251), .Z(n2248) );
  CIVX2 U1480 ( .A(n1985), .Z(n1814) );
  CIVX1 U1481 ( .A(a[24]), .Z(n1993) );
  CIVX2 U1482 ( .A(n2215), .Z(n1978) );
  CNIVX1 U1483 ( .A(n1755), .Z(n1606) );
  CEOX2 U1484 ( .A(n1686), .B(n1683), .Z(n1608) );
  CIVX1 U1485 ( .A(a[22]), .Z(n1833) );
  CIVX1 U1486 ( .A(n1656), .Z(n1657) );
  CNIVX1 U1487 ( .A(n940), .Z(n1609) );
  COR2XL U1488 ( .A(net171503), .B(n481), .Z(n1610) );
  CAN2XL U1489 ( .A(n1543), .B(n873), .Z(n1611) );
  CAN2XL U1490 ( .A(n2007), .B(n332), .Z(product[1]) );
  CENX2 U1491 ( .A(n1969), .B(a[18]), .Z(n1865) );
  COND1X1 U1492 ( .A(n325), .B(n323), .C(n324), .Z(n322) );
  CEOX2 U1493 ( .A(n2194), .B(n544), .Z(n540) );
  COND2X1 U1494 ( .A(n84), .B(n1141), .C(n1864), .D(n1140), .Z(n863) );
  CEOX1 U1495 ( .A(n1889), .B(n863), .Z(n532) );
  CND2XL U1496 ( .A(n992), .B(n946), .Z(n1660) );
  CIVX2 U1497 ( .A(n2243), .Z(n2238) );
  CHA1XL U1498 ( .A(n811), .B(n995), .CO(n785), .S(n786) );
  CND2XL U1499 ( .A(n1948), .B(n1949), .Z(n1613) );
  COND2XL U1500 ( .A(n1147), .B(n2190), .C(n1693), .D(n1146), .Z(n869) );
  COND2X1 U1501 ( .A(n2190), .B(n1145), .C(n1865), .D(n1144), .Z(n867) );
  CND2XL U1502 ( .A(n1412), .B(n1865), .Z(n84) );
  CND2X1 U1503 ( .A(n1412), .B(n1864), .Z(n2190) );
  COR2X1 U1504 ( .A(n512), .B(n535), .Z(n1936) );
  COND2X1 U1505 ( .A(n1905), .B(n1143), .C(n1864), .D(n1142), .Z(n865) );
  CND2XL U1506 ( .A(n681), .B(n670), .Z(n1856) );
  CIVX1 U1507 ( .A(n105), .Z(n1804) );
  CIVXL U1508 ( .A(n1875), .Z(n1614) );
  CENXL U1509 ( .A(n1615), .B(n674), .Z(n672) );
  CND2X1 U1510 ( .A(n1412), .B(n1864), .Z(n1905) );
  CENX1 U1511 ( .A(net33480), .B(n2255), .Z(n1781) );
  CENXL U1512 ( .A(n2201), .B(n2002), .Z(n1180) );
  CFA1XL U1513 ( .A(n858), .B(n948), .CI(n888), .CO(n399), .S(n400) );
  CIVX1 U1514 ( .A(n684), .Z(n1875) );
  CENX1 U1515 ( .A(n425), .B(net171635), .Z(n1685) );
  CENX1 U1516 ( .A(n1685), .B(n1677), .Z(n394) );
  CND2X2 U1517 ( .A(n1745), .B(a[14]), .Z(n1748) );
  CND2X2 U1518 ( .A(n2072), .B(n2059), .Z(n1918) );
  CIVX2 U1519 ( .A(n1432), .Z(net179544) );
  CIVXL U1520 ( .A(n1555), .Z(n1616) );
  CIVX2 U1521 ( .A(n1616), .Z(n1617) );
  CENX1 U1522 ( .A(n2201), .B(n1975), .Z(n1224) );
  CIVXL U1523 ( .A(n61), .Z(n1618) );
  CIVX1 U1524 ( .A(n1618), .Z(n1619) );
  CND2X2 U1525 ( .A(n1415), .B(n58), .Z(n61) );
  CND2X2 U1526 ( .A(n2004), .B(n2005), .Z(n1022) );
  COR2X1 U1527 ( .A(n27), .B(n1307), .Z(n2004) );
  CNR2IX1 U1528 ( .B(net33082), .A(n89), .Z(n856) );
  CFA1X1 U1529 ( .A(n1007), .B(n618), .CI(n635), .CO(n609), .S(n610) );
  CNR2IX2 U1530 ( .B(net33082), .A(n1865), .Z(n870) );
  COND2XL U1531 ( .A(n18), .B(n1320), .C(n1319), .D(n2185), .Z(n1034) );
  COND2XL U1532 ( .A(n18), .B(n1317), .C(n1316), .D(n2185), .Z(n1031) );
  COND2XL U1533 ( .A(n18), .B(n1314), .C(n1313), .D(n2185), .Z(n1028) );
  COND2XL U1534 ( .A(n18), .B(n1316), .C(n1315), .D(n2185), .Z(n1030) );
  COND2XL U1535 ( .A(n18), .B(n1315), .C(n1314), .D(n2185), .Z(n1029) );
  COND2XL U1536 ( .A(n18), .B(n1318), .C(n1317), .D(n2185), .Z(n1032) );
  COND2XL U1537 ( .A(n18), .B(n1323), .C(n1322), .D(n2185), .Z(n1037) );
  COND2XL U1538 ( .A(n18), .B(n1322), .C(n1321), .D(n2185), .Z(n1036) );
  COND2XL U1539 ( .A(n18), .B(n1326), .C(n1325), .D(n2185), .Z(n1040) );
  COND2XL U1540 ( .A(n18), .B(n1329), .C(n1328), .D(n2185), .Z(n1043) );
  CENXL U1541 ( .A(n171), .B(n1620), .Z(product[28]) );
  CAN2XL U1542 ( .A(n336), .B(net179954), .Z(n1620) );
  CIVX2 U1543 ( .A(n2216), .Z(n1771) );
  CIVXL U1544 ( .A(n1834), .Z(n1621) );
  CIVX1 U1545 ( .A(n1963), .Z(n1834) );
  CIVXL U1546 ( .A(n223), .Z(n222) );
  COND2X1 U1547 ( .A(n27), .B(n1305), .C(n1304), .D(n2009), .Z(n1020) );
  CFA1X1 U1548 ( .A(n970), .B(n1020), .CI(n994), .CO(n779), .S(n780) );
  CIVXL U1549 ( .A(n69), .Z(n1622) );
  CIVX2 U1550 ( .A(n1622), .Z(n1623) );
  CND2X2 U1551 ( .A(n1762), .B(n66), .Z(n69) );
  CFA1X1 U1552 ( .A(n1005), .B(n578), .CI(n1033), .CO(n569), .S(n570) );
  CIVX2 U1553 ( .A(n2213), .Z(n1745) );
  CHA1X1 U1554 ( .A(n810), .B(n1077), .CO(n773), .S(n774) );
  CND2XL U1555 ( .A(n104), .B(a[28]), .Z(n1986) );
  CND2XL U1556 ( .A(n682), .B(n693), .Z(n1946) );
  CENXL U1557 ( .A(n1731), .B(n662), .Z(n658) );
  CENX1 U1558 ( .A(n1624), .B(n1579), .Z(n446) );
  CENX1 U1559 ( .A(n2150), .B(n456), .Z(n1624) );
  CENX1 U1560 ( .A(n1625), .B(n1764), .Z(n440) );
  CENXL U1561 ( .A(n446), .B(n469), .Z(n1625) );
  CEOX2 U1562 ( .A(n1636), .B(n447), .Z(n416) );
  COND1X2 U1563 ( .A(n184), .B(n178), .C(n179), .Z(n173) );
  CENX1 U1564 ( .A(n1626), .B(n806), .Z(n684) );
  CENX1 U1565 ( .A(n961), .B(n1069), .Z(n1626) );
  CNIVX4 U1566 ( .A(n71), .Z(n2214) );
  CENX1 U1567 ( .A(n1969), .B(a[18]), .Z(n1864) );
  CND2XL U1568 ( .A(n469), .B(n446), .Z(net180107) );
  CND2X1 U1569 ( .A(n463), .B(n440), .Z(net180482) );
  COND1XL U1570 ( .A(n307), .B(n309), .C(n308), .Z(n1627) );
  COND1X2 U1571 ( .A(n307), .B(n309), .C(n308), .Z(n306) );
  CANR1X2 U1572 ( .A(n314), .B(n2022), .C(n311), .Z(n309) );
  CNIVX1 U1573 ( .A(n1629), .Z(product[12]) );
  CNIVX1 U1574 ( .A(n2258), .Z(n1629) );
  CND2XL U1575 ( .A(n350), .B(n2177), .Z(n136) );
  CNIVX1 U1576 ( .A(n1631), .Z(product[10]) );
  CNIVX1 U1577 ( .A(n2259), .Z(n1631) );
  CND2XL U1578 ( .A(n2028), .B(n252), .Z(n133) );
  CND2XL U1579 ( .A(n2091), .B(n2089), .Z(n252) );
  CIVXL U1580 ( .A(n261), .Z(n260) );
  CNIVXL U1581 ( .A(n2180), .Z(n1632) );
  CND2XL U1582 ( .A(n348), .B(n1632), .Z(n134) );
  CNIVX1 U1583 ( .A(n1634), .Z(product[15]) );
  CNIVX1 U1584 ( .A(n2257), .Z(n1634) );
  CND2XL U1585 ( .A(n2182), .B(n2179), .Z(n135) );
  CIVX3 U1586 ( .A(n2161), .Z(n278) );
  CND2XL U1587 ( .A(n1581), .B(n455), .Z(n1872) );
  CEO3XL U1588 ( .A(n2171), .B(n2069), .C(n2066), .Z(n1699) );
  CND2X1 U1589 ( .A(n2069), .B(n2066), .Z(n1932) );
  CENX2 U1590 ( .A(n1635), .B(n2037), .Z(n480) );
  CENX2 U1591 ( .A(n2079), .B(n2040), .Z(n1635) );
  CND2X1 U1592 ( .A(n498), .B(n519), .Z(n1767) );
  CEOX2 U1593 ( .A(net171634), .B(n449), .Z(n1636) );
  CND2XL U1594 ( .A(n447), .B(n449), .Z(n1637) );
  CND2XL U1595 ( .A(n447), .B(net171634), .Z(n1638) );
  CND2XL U1596 ( .A(n449), .B(net171634), .Z(n1639) );
  CND3XL U1597 ( .A(n1637), .B(n1638), .C(n1639), .Z(n415) );
  CEOX1 U1598 ( .A(n807), .B(n963), .Z(n714) );
  CIVX2 U1599 ( .A(n1640), .Z(n713) );
  CND2X1 U1600 ( .A(n963), .B(n807), .Z(n1640) );
  CENX1 U1601 ( .A(net33482), .B(n2249), .Z(n1251) );
  CNIVX4 U1602 ( .A(n1404), .Z(net33482) );
  COND2X1 U1603 ( .A(n1183), .B(n69), .C(n66), .D(n1182), .Z(n1697) );
  CNR2X1 U1604 ( .A(n167), .B(n162), .Z(n160) );
  CND2X1 U1605 ( .A(n496), .B(n519), .Z(n1768) );
  CEOX2 U1606 ( .A(n1741), .B(n426), .Z(n418) );
  CEOX1 U1607 ( .A(n632), .B(n634), .Z(n1641) );
  CEOXL U1608 ( .A(n1641), .B(n636), .Z(n626) );
  CND2XL U1609 ( .A(n636), .B(n634), .Z(n1642) );
  CND2XL U1610 ( .A(n636), .B(n632), .Z(n1643) );
  CND2X1 U1611 ( .A(n634), .B(n632), .Z(n1644) );
  CND3XL U1612 ( .A(n1642), .B(n1643), .C(n1644), .Z(n625) );
  CENXL U1613 ( .A(net33480), .B(n2215), .Z(n1145) );
  CND2X1 U1614 ( .A(n1942), .B(n1943), .Z(n1408) );
  CEO3XL U1615 ( .A(n899), .B(n805), .C(n869), .Z(n652) );
  CND2X1 U1616 ( .A(n899), .B(n869), .Z(n1645) );
  CEOX1 U1617 ( .A(n649), .B(n647), .Z(n1648) );
  CND2X1 U1618 ( .A(n649), .B(n647), .Z(n1649) );
  CND3XL U1619 ( .A(n1649), .B(n1650), .C(n1651), .Z(n627) );
  CENX2 U1620 ( .A(n1975), .B(n1971), .Z(n1652) );
  CIVX1 U1621 ( .A(n2253), .Z(n2252) );
  CENX2 U1622 ( .A(n1975), .B(n1971), .Z(n58) );
  COND2X1 U1623 ( .A(n77), .B(n1161), .C(n74), .D(n1160), .Z(n882) );
  CND2X1 U1624 ( .A(n1545), .B(n456), .Z(n1653) );
  CND2X1 U1625 ( .A(n456), .B(n2150), .Z(n1655) );
  CND3X2 U1626 ( .A(n1653), .B(n1654), .C(n1655), .Z(n445) );
  CND2XL U1627 ( .A(n921), .B(n1071), .Z(n1883) );
  CND2X1 U1628 ( .A(n1410), .B(n95), .Z(n1669) );
  CENX1 U1629 ( .A(n664), .B(n675), .Z(n1731) );
  CIVX1 U1630 ( .A(n301), .Z(n300) );
  CANR1X2 U1631 ( .A(n2018), .B(n306), .C(n303), .Z(n301) );
  CIVXL U1632 ( .A(n1965), .Z(n1722) );
  CIVX3 U1633 ( .A(n1965), .Z(n1971) );
  CND2IX1 U1634 ( .B(a[18]), .A(n2215), .Z(n1980) );
  CENX1 U1635 ( .A(n479), .B(n2149), .Z(n1851) );
  CND3X1 U1636 ( .A(n1997), .B(n1998), .C(n1999), .Z(n1658) );
  CND2X1 U1637 ( .A(n2170), .B(n2065), .Z(n1997) );
  CND2XL U1638 ( .A(n968), .B(n992), .Z(n1659) );
  CND2XL U1639 ( .A(n968), .B(n946), .Z(n1661) );
  CND3XL U1640 ( .A(n1659), .B(n1660), .C(n1661), .Z(n765) );
  CANR1X1 U1641 ( .A(n297), .B(n2014), .C(n292), .Z(n1966) );
  CND2X1 U1642 ( .A(n2014), .B(n2016), .Z(n289) );
  CND3X1 U1643 ( .A(n1997), .B(n1998), .C(n1999), .Z(n509) );
  CND2X1 U1644 ( .A(n2170), .B(n2068), .Z(n1998) );
  CAN2X1 U1645 ( .A(n223), .B(n187), .Z(n1939) );
  CNR2XL U1646 ( .A(n1597), .B(n1937), .Z(n1662) );
  CIVX2 U1647 ( .A(n294), .Z(n292) );
  CIVXL U1648 ( .A(n184), .Z(n182) );
  CENXL U1649 ( .A(n185), .B(n124), .Z(product[26]) );
  CENX2 U1650 ( .A(n529), .B(n1663), .Z(n500) );
  CENX1 U1651 ( .A(n527), .B(n2138), .Z(n1663) );
  CEOX1 U1652 ( .A(n2125), .B(n2124), .Z(n1664) );
  CEOX1 U1653 ( .A(n1664), .B(n574), .Z(n566) );
  CND2XL U1654 ( .A(n574), .B(n2124), .Z(n1665) );
  CND2XL U1655 ( .A(n574), .B(n2125), .Z(n1666) );
  CND2XL U1656 ( .A(n2124), .B(n2125), .Z(n1667) );
  CND3X2 U1657 ( .A(n1665), .B(n1666), .C(n1667), .Z(n565) );
  CENX1 U1658 ( .A(n2052), .B(n1866), .Z(n574) );
  CEOX2 U1659 ( .A(n546), .B(n565), .Z(n2194) );
  CENX1 U1660 ( .A(n2070), .B(n2049), .Z(n1866) );
  CIVX2 U1661 ( .A(n104), .Z(n1985) );
  CND2XL U1662 ( .A(n816), .B(n846), .Z(n1951) );
  CENXL U1663 ( .A(n2205), .B(n2217), .Z(n1668) );
  CNIVX4 U1664 ( .A(n1402), .Z(n2201) );
  CENX1 U1665 ( .A(n2240), .B(n2201), .Z(n1276) );
  CENXL U1666 ( .A(n2233), .B(n2201), .Z(n1305) );
  CENXL U1667 ( .A(n2247), .B(n2201), .Z(n1249) );
  COND2XL U1668 ( .A(n61), .B(n1202), .C(n1652), .D(n1201), .Z(n921) );
  CEOX1 U1669 ( .A(n2143), .B(n2140), .Z(n1670) );
  CND2X1 U1670 ( .A(n510), .B(n2140), .Z(n1671) );
  CND2X1 U1671 ( .A(n510), .B(n2143), .Z(n1672) );
  CND2XL U1672 ( .A(n2140), .B(n2143), .Z(n1673) );
  CND3X2 U1673 ( .A(n1671), .B(n1672), .C(n1673), .Z(n497) );
  COND2XL U1674 ( .A(n1669), .B(n1668), .C(n95), .D(n1111), .Z(n1674) );
  CNIVX2 U1675 ( .A(n93), .Z(n2217) );
  CND2IX2 U1676 ( .B(n2006), .A(n74), .Z(n77) );
  CIVXL U1677 ( .A(n1964), .Z(n1675) );
  CIVX2 U1678 ( .A(n1675), .Z(n1676) );
  CENX1 U1679 ( .A(net33480), .B(n1975), .Z(n1225) );
  CND2XL U1680 ( .A(n941), .B(n1071), .Z(n1884) );
  CND2XL U1681 ( .A(n941), .B(n921), .Z(n1882) );
  CIVX8 U1682 ( .A(n2256), .Z(n2254) );
  CND2X1 U1683 ( .A(n2065), .B(n2068), .Z(n1999) );
  COND1X2 U1684 ( .A(n1678), .B(n1679), .C(n1680), .Z(n1677) );
  CNR2X2 U1685 ( .A(n1681), .B(n1682), .Z(n393) );
  CIVX2 U1686 ( .A(net171723), .Z(n1683) );
  CIVX2 U1687 ( .A(net171759), .Z(n1678) );
  CIVX2 U1688 ( .A(n425), .Z(n1684) );
  CENX2 U1689 ( .A(net182724), .B(n1608), .Z(n420) );
  CENX2 U1690 ( .A(net171738), .B(net171759), .Z(n1686) );
  CIVX2 U1691 ( .A(n1688), .Z(n1687) );
  CIVXL U1692 ( .A(net171738), .Z(n1688) );
  COND1X1 U1693 ( .A(n1690), .B(net179954), .C(n163), .Z(n1689) );
  CANR1X1 U1694 ( .A(n173), .B(net179971), .C(n1689), .Z(net179515) );
  COND1XL U1695 ( .A(net179954), .B(n1690), .C(n163), .Z(net180013) );
  CND2X2 U1696 ( .A(n408), .B(n435), .Z(n163) );
  CAN2XL U1697 ( .A(n163), .B(n335), .Z(net179680) );
  CND2X1 U1698 ( .A(n380), .B(n407), .Z(n156) );
  COR2X1 U1699 ( .A(n407), .B(n380), .Z(net178620) );
  CND2X2 U1700 ( .A(net182663), .B(net182662), .Z(n422) );
  CND3X1 U1701 ( .A(net180105), .B(net180106), .C(net180107), .Z(n439) );
  CNIVX2 U1702 ( .A(n412), .Z(net179910) );
  CEOXL U1703 ( .A(n1691), .B(n438), .Z(n436) );
  CEOXL U1704 ( .A(n440), .B(n463), .Z(n1691) );
  CND2X2 U1705 ( .A(n462), .B(n487), .Z(n179) );
  CND2X1 U1706 ( .A(n438), .B(n463), .Z(net180480) );
  CEO3X1 U1707 ( .A(n440), .B(net179996), .C(n1551), .Z(net179805) );
  CNR2X2 U1708 ( .A(net179493), .B(n435), .Z(n162) );
  CANR1X1 U1709 ( .A(net178620), .B(net179430), .C(n154), .Z(n152) );
  CENXL U1710 ( .A(net179380), .B(n152), .Z(product[31]) );
  CND2X1 U1711 ( .A(net179515), .B(net179197), .Z(net179430) );
  CIVX2 U1712 ( .A(n173), .Z(n175) );
  COND1XL U1713 ( .A(n167), .B(n175), .C(net179954), .Z(n166) );
  CNR2X1 U1714 ( .A(net179834), .B(n487), .Z(n178) );
  COR2X1 U1715 ( .A(n158), .B(n186), .Z(net179197) );
  CND2XL U1716 ( .A(n159), .B(net179197), .Z(n157) );
  CND2X1 U1717 ( .A(n160), .B(n172), .Z(n158) );
  CNR2XL U1718 ( .A(n167), .B(n162), .Z(net179971) );
  CANR1XL U1719 ( .A(n173), .B(net179971), .C(net180013), .Z(n159) );
  CND2XL U1720 ( .A(net171639), .B(net171637), .Z(net180018) );
  CND2XL U1721 ( .A(n1608), .B(net171637), .Z(net180017) );
  CND2XL U1722 ( .A(n1608), .B(net171639), .Z(net180016) );
  CNIVX1 U1723 ( .A(n1865), .Z(n1693) );
  CENX1 U1724 ( .A(a[6]), .B(n2245), .Z(n1418) );
  CIVX2 U1725 ( .A(n30), .Z(n2245) );
  CND2XL U1726 ( .A(n566), .B(n564), .Z(n1728) );
  CND3X2 U1727 ( .A(n1920), .B(n1919), .C(n1918), .Z(n505) );
  CNIVX1 U1728 ( .A(n79), .Z(n1694) );
  CNIVX4 U1729 ( .A(n79), .Z(n2215) );
  CIVXL U1730 ( .A(n530), .Z(n1695) );
  CIVXL U1731 ( .A(n1695), .Z(n1696) );
  CFA1XL U1732 ( .A(n862), .B(n930), .CI(n876), .CO(n507), .S(n508) );
  CIVXL U1733 ( .A(n1561), .Z(n1698) );
  CND3X1 U1734 ( .A(n2198), .B(n2199), .C(n2200), .Z(n535) );
  CENX1 U1735 ( .A(n1769), .B(n514), .Z(n512) );
  CENX1 U1736 ( .A(n537), .B(n516), .Z(n1769) );
  CND2X2 U1737 ( .A(n1702), .B(n1703), .Z(n1783) );
  CIVX1 U1738 ( .A(n2068), .Z(n1700) );
  CIVX2 U1739 ( .A(n2065), .Z(n1701) );
  CND2IX4 U1740 ( .B(n2008), .A(n2009), .Z(n27) );
  COND2X1 U1741 ( .A(n27), .B(n1303), .C(n1302), .D(n2009), .Z(n1018) );
  CEO3X2 U1742 ( .A(n2162), .B(n2114), .C(n2112), .Z(n590) );
  CND2X1 U1743 ( .A(n2162), .B(n2114), .Z(n1704) );
  CND2X1 U1744 ( .A(n2162), .B(n2112), .Z(n1705) );
  CND2X1 U1745 ( .A(n2114), .B(n2112), .Z(n1706) );
  CND3X2 U1746 ( .A(n1704), .B(n1705), .C(n1706), .Z(n589) );
  CEOX2 U1747 ( .A(n2126), .B(n2128), .Z(n1707) );
  CEOX2 U1748 ( .A(n1707), .B(n589), .Z(n564) );
  CND2XL U1749 ( .A(n2126), .B(n2128), .Z(n1708) );
  CND2XL U1750 ( .A(n2126), .B(n589), .Z(n1709) );
  CND2XL U1751 ( .A(n2128), .B(n589), .Z(n1710) );
  CND3X1 U1752 ( .A(n1708), .B(n1709), .C(n1710), .Z(n563) );
  CND2X1 U1753 ( .A(n1761), .B(n583), .Z(n1713) );
  CND2X2 U1754 ( .A(n1711), .B(n1712), .Z(n1714) );
  CND2X2 U1755 ( .A(n1713), .B(n1714), .Z(n560) );
  CIVX2 U1756 ( .A(n1761), .Z(n1711) );
  CIVXL U1757 ( .A(n583), .Z(n1712) );
  CND2X1 U1758 ( .A(n1696), .B(n528), .Z(n1897) );
  COND2XL U1759 ( .A(n44), .B(n1238), .C(n1237), .D(n42), .Z(n955) );
  COND2XL U1760 ( .A(n44), .B(n1230), .C(n1229), .D(n42), .Z(n947) );
  COND2XL U1761 ( .A(n44), .B(n1232), .C(n1231), .D(n42), .Z(n949) );
  COND2XL U1762 ( .A(n44), .B(n1240), .C(n1239), .D(n42), .Z(n957) );
  COND2XL U1763 ( .A(n44), .B(n1231), .C(n1230), .D(n42), .Z(n948) );
  COND2XL U1764 ( .A(n44), .B(n1239), .C(n1238), .D(n42), .Z(n956) );
  COND2XL U1765 ( .A(n44), .B(n1233), .C(n1232), .D(n42), .Z(n950) );
  COND2XL U1766 ( .A(n44), .B(n1241), .C(n1240), .D(n42), .Z(n958) );
  COND2XL U1767 ( .A(n44), .B(n1235), .C(n1234), .D(n42), .Z(n952) );
  COND2XL U1768 ( .A(n44), .B(n1237), .C(n1236), .D(n42), .Z(n954) );
  COND2XL U1769 ( .A(n44), .B(n1242), .C(n1241), .D(n42), .Z(n959) );
  COND2XL U1770 ( .A(n44), .B(n1243), .C(n1242), .D(n42), .Z(n960) );
  COND2XL U1771 ( .A(n44), .B(n1245), .C(n1244), .D(n42), .Z(n962) );
  COND2XL U1772 ( .A(n44), .B(n1246), .C(n1245), .D(n42), .Z(n963) );
  COND2XL U1773 ( .A(n44), .B(n1247), .C(n1246), .D(n42), .Z(n964) );
  COND2XL U1774 ( .A(n44), .B(n1249), .C(n1248), .D(n42), .Z(n966) );
  COND2XL U1775 ( .A(n44), .B(n1248), .C(n1247), .D(n42), .Z(n965) );
  CIVX1 U1776 ( .A(n299), .Z(n297) );
  CIVX8 U1777 ( .A(n2237), .Z(n2234) );
  CEOX1 U1778 ( .A(n2145), .B(n2147), .Z(n1715) );
  CEOX2 U1779 ( .A(n1715), .B(n506), .Z(n496) );
  CND2XL U1780 ( .A(n506), .B(n2147), .Z(n1716) );
  CND2XL U1781 ( .A(n506), .B(n2145), .Z(n1717) );
  CND2XL U1782 ( .A(n2147), .B(n2145), .Z(n1718) );
  CNIVX2 U1783 ( .A(n63), .Z(n2213) );
  CEOXL U1784 ( .A(n2186), .B(n1035), .Z(n612) );
  CND3X1 U1785 ( .A(n1719), .B(n1720), .C(n1721), .Z(n457) );
  CENX1 U1786 ( .A(n459), .B(n457), .Z(n1780) );
  CENXL U1787 ( .A(n2240), .B(n2202), .Z(n1275) );
  CIVX4 U1788 ( .A(n2244), .Z(n2240) );
  CND2X1 U1789 ( .A(n1965), .B(n2254), .Z(n1724) );
  CND2X2 U1790 ( .A(n1722), .B(n1723), .Z(n1725) );
  CND2X2 U1791 ( .A(n1724), .B(n1725), .Z(n1415) );
  CIVX2 U1792 ( .A(n2254), .Z(n1723) );
  CENXL U1793 ( .A(n2206), .B(n2217), .Z(n1111) );
  CENXL U1794 ( .A(n1963), .B(net33480), .Z(n1117) );
  CENXL U1795 ( .A(n2205), .B(n2217), .Z(n1112) );
  CIVX1 U1796 ( .A(n566), .Z(n1726) );
  CIVX2 U1797 ( .A(n564), .Z(n1727) );
  CENX2 U1798 ( .A(n1730), .B(n2063), .Z(n456) );
  CENX2 U1799 ( .A(n2080), .B(n2056), .Z(n1730) );
  CENX1 U1800 ( .A(n2072), .B(n1782), .Z(n506) );
  CND2X1 U1801 ( .A(a[22]), .B(n1834), .Z(n1835) );
  COND2X1 U1802 ( .A(n44), .B(n1251), .C(n42), .D(n1250), .Z(n968) );
  CNR2IX2 U1803 ( .B(net33082), .A(n100), .Z(n834) );
  CND2XL U1804 ( .A(n806), .B(n1069), .Z(n1852) );
  CND2XL U1805 ( .A(n806), .B(n961), .Z(n1853) );
  CENXL U1806 ( .A(n2220), .B(b[31]), .Z(n1341) );
  CENXL U1807 ( .A(n2220), .B(n1387), .Z(n1354) );
  CENXL U1808 ( .A(n2220), .B(n2203), .Z(n1367) );
  CENXL U1809 ( .A(n2220), .B(n2202), .Z(n1368) );
  CENXL U1810 ( .A(n2220), .B(n2204), .Z(n1366) );
  CENXL U1811 ( .A(n2220), .B(n2201), .Z(n1369) );
  CENXL U1812 ( .A(n2220), .B(net33480), .Z(n1370) );
  CENXL U1813 ( .A(n2220), .B(net33482), .Z(n1371) );
  CENXL U1814 ( .A(n2220), .B(n2206), .Z(n1364) );
  CENXL U1815 ( .A(n2220), .B(n1396), .Z(n1363) );
  CENXL U1816 ( .A(n2220), .B(n2207), .Z(n1362) );
  CENXL U1817 ( .A(n2220), .B(n2208), .Z(n1361) );
  CEOX4 U1818 ( .A(n2220), .B(a[2]), .Z(n2033) );
  CIVX3 U1819 ( .A(n2222), .Z(n2221) );
  CND2X1 U1820 ( .A(n438), .B(n440), .Z(n1843) );
  CND2X1 U1821 ( .A(n498), .B(n496), .Z(n1766) );
  CENX1 U1822 ( .A(n2054), .B(n2059), .Z(n1782) );
  COND2X1 U1823 ( .A(n69), .B(n1181), .C(n1607), .D(n1180), .Z(n901) );
  CENXL U1824 ( .A(n2207), .B(n1698), .Z(n1173) );
  CENXL U1825 ( .A(n2206), .B(n1698), .Z(n1175) );
  CENXL U1826 ( .A(n2211), .B(n1698), .Z(n1169) );
  CENXL U1827 ( .A(n2204), .B(n1560), .Z(n1177) );
  CEOX2 U1828 ( .A(n870), .B(n900), .Z(n1732) );
  CEOX2 U1829 ( .A(n1732), .B(n884), .Z(n670) );
  CND2XL U1830 ( .A(n884), .B(n870), .Z(n1733) );
  CND2XL U1831 ( .A(n884), .B(n900), .Z(n1734) );
  CND2XL U1832 ( .A(n870), .B(n900), .Z(n1735) );
  CND3X1 U1833 ( .A(n1733), .B(n1734), .C(n1735), .Z(n669) );
  CND2X1 U1834 ( .A(n1862), .B(n1863), .Z(n884) );
  CENX1 U1835 ( .A(n476), .B(n1736), .Z(n468) );
  CENX1 U1836 ( .A(n497), .B(n474), .Z(n1736) );
  CND2IX2 U1837 ( .B(n455), .A(n1765), .Z(net182663) );
  CND2XL U1838 ( .A(net182662), .B(net182663), .Z(net184228) );
  CENX4 U1839 ( .A(n2244), .B(a[8]), .Z(n2032) );
  CND2X1 U1840 ( .A(n2062), .B(n2073), .Z(n1738) );
  CND2X1 U1841 ( .A(n2062), .B(n2055), .Z(n1739) );
  CND2X1 U1842 ( .A(n2073), .B(n2055), .Z(n1740) );
  CND3X2 U1843 ( .A(n1738), .B(n1739), .C(n1740), .Z(n481) );
  CND3X1 U1844 ( .A(n1742), .B(n1743), .C(n1744), .Z(n417) );
  CND2X1 U1845 ( .A(n2213), .B(n1746), .Z(n1747) );
  CND2X2 U1846 ( .A(n1747), .B(n1748), .Z(n1762) );
  CIVXL U1847 ( .A(a[14]), .Z(n1746) );
  CND3X2 U1848 ( .A(n1749), .B(n1750), .C(n1751), .Z(n479) );
  CIVX2 U1849 ( .A(a[12]), .Z(n1965) );
  CNIVX4 U1850 ( .A(n79), .Z(n1752) );
  CIVXL U1851 ( .A(n457), .Z(n1753) );
  CIVXL U1852 ( .A(n1753), .Z(n1754) );
  CNIVX4 U1853 ( .A(n86), .Z(n1755) );
  CENXL U1854 ( .A(n2201), .B(n1694), .Z(n1144) );
  CND2X1 U1855 ( .A(n1990), .B(n1991), .Z(n902) );
  CENX2 U1856 ( .A(n2067), .B(n1756), .Z(n530) );
  CND2X1 U1857 ( .A(n1800), .B(n1796), .Z(n1759) );
  CND2X2 U1858 ( .A(n1757), .B(n1758), .Z(n1760) );
  CND2X2 U1859 ( .A(n1759), .B(n1760), .Z(n450) );
  CIVX1 U1860 ( .A(n1800), .Z(n1757) );
  CIVXL U1861 ( .A(n1796), .Z(n1758) );
  CENX1 U1862 ( .A(net171503), .B(n481), .Z(n1800) );
  CENX1 U1863 ( .A(net33482), .B(n1969), .Z(n1163) );
  CNIVX3 U1864 ( .A(n116), .Z(net33080) );
  CENXL U1865 ( .A(net33080), .B(n2249), .Z(n1252) );
  CNR2X2 U1866 ( .A(n750), .B(n759), .Z(n285) );
  CIVXL U1867 ( .A(n467), .Z(n1763) );
  CIVX1 U1868 ( .A(n1763), .Z(n1764) );
  COR2XL U1869 ( .A(n69), .B(n1182), .Z(n1990) );
  CND2X1 U1870 ( .A(n1780), .B(n455), .Z(net182662) );
  CEO3X2 U1871 ( .A(n498), .B(n519), .C(n496), .Z(n492) );
  CND3X2 U1872 ( .A(n1766), .B(n1767), .C(n1768), .Z(n491) );
  CEO3X1 U1873 ( .A(n470), .B(n491), .C(net180095), .Z(n1960) );
  CEOXL U1874 ( .A(net33080), .B(n2253), .Z(n1227) );
  CHA1X1 U1875 ( .A(n945), .B(n809), .CO(n757), .S(n758) );
  COND2X1 U1876 ( .A(n53), .B(n2253), .C(n50), .D(n1228), .Z(n809) );
  CIVX3 U1877 ( .A(n48), .Z(n2253) );
  CENX1 U1878 ( .A(net33080), .B(n2002), .Z(n1183) );
  CND2X2 U1879 ( .A(n1771), .B(a[20]), .Z(n1772) );
  CND2X2 U1880 ( .A(n1755), .B(n1770), .Z(n1773) );
  CIVX2 U1881 ( .A(a[20]), .Z(n1770) );
  COND2XL U1882 ( .A(n1087), .B(n115), .C(n1558), .D(n1086), .Z(n815) );
  CENXL U1883 ( .A(net33080), .B(n113), .Z(n1087) );
  COND2XL U1884 ( .A(n1558), .B(n1088), .C(n1431), .D(n115), .Z(n799) );
  CND2X2 U1885 ( .A(n1432), .B(n1775), .Z(n1777) );
  CIVX2 U1886 ( .A(a[30]), .Z(n1775) );
  CND2X1 U1887 ( .A(n109), .B(a[30]), .Z(n1776) );
  CND2IXL U1888 ( .B(net33082), .A(n113), .Z(n1088) );
  CIVXL U1889 ( .A(n113), .Z(n1431) );
  CENXL U1890 ( .A(net33480), .B(n109), .Z(n1090) );
  CIVXL U1891 ( .A(n1940), .Z(n1778) );
  CND2X1 U1892 ( .A(n488), .B(n511), .Z(n184) );
  CIVX3 U1893 ( .A(n2256), .Z(n2255) );
  CANR1XL U1894 ( .A(n165), .B(n185), .C(n166), .Z(n164) );
  CND2X1 U1895 ( .A(n693), .B(n1875), .Z(n1876) );
  CND2XL U1896 ( .A(n1988), .B(n1989), .Z(n1984) );
  CNR2X2 U1897 ( .A(n91), .B(n1124), .Z(n2000) );
  CENX1 U1898 ( .A(n2206), .B(n2216), .Z(n1124) );
  CENX1 U1899 ( .A(n2203), .B(n1975), .Z(n1222) );
  CEOX1 U1900 ( .A(n933), .B(n879), .Z(n1784) );
  CEOXL U1901 ( .A(n853), .B(n1784), .Z(n576) );
  CND2X1 U1902 ( .A(n853), .B(n879), .Z(n1785) );
  CND2X1 U1903 ( .A(n853), .B(n933), .Z(n1786) );
  CND2X1 U1904 ( .A(n879), .B(n933), .Z(n1787) );
  CND3X2 U1905 ( .A(n1785), .B(n1786), .C(n1787), .Z(n575) );
  CNR2X2 U1906 ( .A(n1789), .B(n1788), .Z(n471) );
  CNR2IX2 U1907 ( .B(n1610), .A(n1790), .Z(n449) );
  CIVX2 U1908 ( .A(net171725), .Z(n1791) );
  CIVX2 U1909 ( .A(net171708), .Z(n1792) );
  CIVX2 U1910 ( .A(net171643), .Z(n1793) );
  CNR2IX2 U1911 ( .B(n1793), .A(n1794), .Z(n1788) );
  CANR1X2 U1912 ( .A(net171643), .B(n1794), .C(n480), .Z(n1789) );
  CNR2X2 U1913 ( .A(net171725), .B(net171752), .Z(n1795) );
  COND1X2 U1914 ( .A(n1792), .B(n1795), .C(n1797), .Z(n1796) );
  CENX2 U1915 ( .A(n1799), .B(n1791), .Z(n1798) );
  CND2X2 U1916 ( .A(net171725), .B(net171752), .Z(n1797) );
  CIVX2 U1917 ( .A(n1798), .Z(n1794) );
  CENX2 U1918 ( .A(net171752), .B(net171708), .Z(n1799) );
  CAN2XL U1919 ( .A(n481), .B(net171503), .Z(n1801) );
  CNR2X2 U1920 ( .A(n1801), .B(n1796), .Z(n1790) );
  CND2X1 U1921 ( .A(n379), .B(n364), .Z(n151) );
  COR2X1 U1922 ( .A(n379), .B(n364), .Z(n1802) );
  CEO3X2 U1923 ( .A(n412), .B(n1803), .C(n437), .Z(net179493) );
  CEO3X1 U1924 ( .A(n1779), .B(net179947), .C(net179913), .Z(n1803) );
  COND2X1 U1925 ( .A(n61), .B(n1781), .C(n1652), .D(n1201), .Z(n1806) );
  CND2XL U1926 ( .A(n1986), .B(n1987), .Z(n1807) );
  CENX1 U1927 ( .A(a[8]), .B(n2250), .Z(n1417) );
  CEOXL U1928 ( .A(net33482), .B(n2253), .Z(n1226) );
  CENXL U1929 ( .A(net33482), .B(n1963), .Z(n1118) );
  COND2X1 U1930 ( .A(n61), .B(n1203), .C(n1652), .D(n1781), .Z(n922) );
  CEO3X2 U1931 ( .A(n2084), .B(n2048), .C(n2046), .Z(n426) );
  CND2XL U1932 ( .A(n2084), .B(n2046), .Z(n1808) );
  CND2XL U1933 ( .A(n2084), .B(n2048), .Z(n1809) );
  CND2X1 U1934 ( .A(n2046), .B(n2048), .Z(n1810) );
  CND3X1 U1935 ( .A(n1808), .B(n1809), .C(n1810), .Z(n425) );
  CNR2IX1 U1936 ( .B(net33082), .A(n66), .Z(n904) );
  CND2XL U1937 ( .A(n843), .B(n979), .Z(n1811) );
  CND2XL U1938 ( .A(n843), .B(n1063), .Z(n1812) );
  CND2X1 U1939 ( .A(n979), .B(n1063), .Z(n1813) );
  CND3XL U1940 ( .A(n1811), .B(n1812), .C(n1813), .Z(n571) );
  COND2XL U1941 ( .A(n9), .B(n1350), .C(n6), .D(n1349), .Z(n1063) );
  COND2XL U1942 ( .A(n1669), .B(n1119), .C(n95), .D(n1118), .Z(n843) );
  COND2XL U1943 ( .A(n1107), .B(n102), .C(n1984), .D(n1106), .Z(n832) );
  CNR2XL U1944 ( .A(n740), .B(n749), .Z(n1815) );
  CNR2XL U1945 ( .A(n740), .B(n749), .Z(n282) );
  CENXL U1946 ( .A(n2252), .B(n2208), .Z(n1216) );
  CENXL U1947 ( .A(n2252), .B(n2207), .Z(n1217) );
  CENXL U1948 ( .A(n2252), .B(n2206), .Z(n1219) );
  CENXL U1949 ( .A(n2252), .B(n1396), .Z(n1218) );
  CENXL U1950 ( .A(n2252), .B(n2209), .Z(n1215) );
  CENXL U1951 ( .A(n2252), .B(n2210), .Z(n1214) );
  CENXL U1952 ( .A(n2252), .B(n2212), .Z(n1212) );
  CENXL U1953 ( .A(n2252), .B(n2211), .Z(n1213) );
  CENXL U1954 ( .A(n2252), .B(n1389), .Z(n1211) );
  CENXL U1955 ( .A(n2252), .B(n1388), .Z(n1210) );
  CIVX1 U1956 ( .A(n2218), .Z(n1994) );
  COND2XL U1957 ( .A(n1183), .B(n69), .C(n1607), .D(n1182), .Z(n1816) );
  CND2X1 U1958 ( .A(n2078), .B(n2053), .Z(n1959) );
  CND3X2 U1959 ( .A(n1957), .B(n1958), .C(n1959), .Z(n529) );
  CND2X1 U1960 ( .A(n2067), .B(n2053), .Z(n1958) );
  CIVX1 U1961 ( .A(net180094), .Z(net180095) );
  CEO3X2 U1962 ( .A(n680), .B(n691), .C(n678), .Z(n674) );
  CND2XL U1963 ( .A(n680), .B(n691), .Z(n1817) );
  CND2XL U1964 ( .A(n680), .B(n678), .Z(n1818) );
  CND2X1 U1965 ( .A(n691), .B(n678), .Z(n1819) );
  CND3XL U1966 ( .A(n1817), .B(n1818), .C(n1819), .Z(n673) );
  CND2XL U1967 ( .A(n689), .B(n676), .Z(n1820) );
  CND2XL U1968 ( .A(n689), .B(n674), .Z(n1821) );
  CND2XL U1969 ( .A(n676), .B(n674), .Z(n1822) );
  CND3XL U1970 ( .A(n1820), .B(n1821), .C(n1822), .Z(n671) );
  CENXL U1971 ( .A(n2242), .B(n1388), .Z(n1262) );
  CENXL U1972 ( .A(n2242), .B(n1387), .Z(n1261) );
  CENXL U1973 ( .A(net33080), .B(n2242), .Z(n1279) );
  CIVX2 U1974 ( .A(n2245), .Z(n2242) );
  COND2X1 U1975 ( .A(n1109), .B(n1984), .C(n1994), .D(n102), .Z(n802) );
  CENX2 U1976 ( .A(n2139), .B(n530), .Z(n1823) );
  CND2X1 U1977 ( .A(n1992), .B(n2170), .Z(n1825) );
  CND2X2 U1978 ( .A(n1783), .B(n1824), .Z(n1826) );
  CND2X2 U1979 ( .A(n1825), .B(n1826), .Z(n510) );
  CIVXL U1980 ( .A(n2170), .Z(n1824) );
  CND2XL U1981 ( .A(n514), .B(n516), .Z(n1827) );
  CND2XL U1982 ( .A(n514), .B(n537), .Z(n1828) );
  CND2XL U1983 ( .A(n516), .B(n537), .Z(n1829) );
  CND3XL U1984 ( .A(n1827), .B(n1828), .C(n1829), .Z(n511) );
  CEO3X1 U1985 ( .A(n2133), .B(n2163), .C(n2131), .Z(n524) );
  CND2X1 U1986 ( .A(n2133), .B(n2131), .Z(n1830) );
  CND2X1 U1987 ( .A(n2133), .B(n2163), .Z(n1831) );
  CND2X1 U1988 ( .A(n2131), .B(n2163), .Z(n1832) );
  CND3X2 U1989 ( .A(n1830), .B(n1831), .C(n1832), .Z(n523) );
  CENX1 U1990 ( .A(n2137), .B(n524), .Z(n1867) );
  CND2XL U1991 ( .A(n1755), .B(a[22]), .Z(n1973) );
  CND2X1 U1992 ( .A(n1963), .B(n1833), .Z(n1836) );
  CND2X2 U1993 ( .A(n1835), .B(n1836), .Z(n1410) );
  CND2X1 U1994 ( .A(n2035), .B(n1658), .Z(n1837) );
  CND2X1 U1995 ( .A(n1658), .B(n2164), .Z(n1839) );
  CND2XL U1996 ( .A(n474), .B(n497), .Z(n1840) );
  CND2XL U1997 ( .A(n474), .B(n476), .Z(n1841) );
  CND2XL U1998 ( .A(n497), .B(n476), .Z(n1842) );
  CND3X1 U1999 ( .A(n1840), .B(n1841), .C(n1842), .Z(n467) );
  CND3X2 U2000 ( .A(net180480), .B(n1843), .C(net180482), .Z(n435) );
  CND3XL U2001 ( .A(net180105), .B(net180106), .C(net180107), .Z(net180475) );
  CND2X4 U2002 ( .A(n1416), .B(n50), .Z(n53) );
  CIVXL U2003 ( .A(n285), .Z(n353) );
  COND2X1 U2004 ( .A(n18), .B(n1332), .C(n1331), .D(n2185), .Z(n1046) );
  COR2X1 U2005 ( .A(n558), .B(n579), .Z(n1844) );
  CEO3X2 U2006 ( .A(n607), .B(n605), .C(n590), .Z(n584) );
  CND2X1 U2007 ( .A(n607), .B(n590), .Z(n1846) );
  CND3X2 U2008 ( .A(n1845), .B(n1846), .C(n1847), .Z(n583) );
  CND2XL U2009 ( .A(n566), .B(n564), .Z(n1848) );
  CND2XL U2010 ( .A(n566), .B(n583), .Z(n1849) );
  CND2XL U2011 ( .A(n564), .B(n583), .Z(n1850) );
  CND3X1 U2012 ( .A(n1848), .B(n1849), .C(n1850), .Z(n559) );
  CND2XL U2013 ( .A(n337), .B(n179), .Z(n123) );
  CENX1 U2014 ( .A(net33482), .B(n1694), .Z(n1146) );
  CIVX1 U2015 ( .A(a[28]), .Z(net179371) );
  CENX2 U2016 ( .A(a[10]), .B(n2253), .Z(n1416) );
  CND2X1 U2017 ( .A(n544), .B(n546), .Z(n2196) );
  CND2XL U2018 ( .A(n1069), .B(n961), .Z(n1854) );
  COND2XL U2019 ( .A(n9), .B(n1356), .C(n6), .D(n1355), .Z(n1069) );
  COND2XL U2020 ( .A(n44), .B(n1244), .C(n1243), .D(n42), .Z(n961) );
  CND2XL U2021 ( .A(n1874), .B(n684), .Z(n1877) );
  CEOXL U2022 ( .A(n1899), .B(n1816), .Z(n710) );
  COR2XL U2023 ( .A(n1607), .B(n1181), .Z(n1991) );
  COND2X1 U2024 ( .A(n61), .B(n2256), .C(n58), .D(n1205), .Z(n808) );
  CEOX2 U2025 ( .A(n2218), .B(n1940), .Z(n105) );
  CIVX1 U2026 ( .A(a[26]), .Z(n1940) );
  CENXL U2027 ( .A(n2003), .B(n1855), .Z(product[11]) );
  CAN2X1 U2028 ( .A(n353), .B(n286), .Z(n1855) );
  CHA1X1 U2029 ( .A(n901), .B(n939), .CO(n685), .S(n686) );
  COND2X1 U2030 ( .A(n1227), .B(n53), .C(n50), .D(n1226), .Z(n945) );
  CEO3X2 U2031 ( .A(n681), .B(n670), .C(n668), .Z(n662) );
  CND2XL U2032 ( .A(n681), .B(n668), .Z(n1857) );
  CND2X1 U2033 ( .A(n670), .B(n668), .Z(n1858) );
  CND3X1 U2034 ( .A(n1856), .B(n1857), .C(n1858), .Z(n661) );
  CND2XL U2035 ( .A(n664), .B(n675), .Z(n1859) );
  CND2XL U2036 ( .A(n664), .B(n662), .Z(n1860) );
  CND2XL U2037 ( .A(n675), .B(n662), .Z(n1861) );
  CND3XL U2038 ( .A(n1859), .B(n1860), .C(n1861), .Z(n657) );
  COR2X1 U2039 ( .A(n77), .B(n1163), .Z(n1862) );
  COR2X1 U2040 ( .A(n74), .B(n1162), .Z(n1863) );
  CENX2 U2041 ( .A(n1560), .B(a[16]), .Z(n74) );
  CENXL U2042 ( .A(net33480), .B(n1969), .Z(n1162) );
  CFA1XL U2043 ( .A(n1021), .B(n1079), .CI(n1049), .CO(n783), .S(n784) );
  COND2X1 U2044 ( .A(n18), .B(n1335), .C(n1334), .D(n2185), .Z(n1049) );
  CFA1XL U2045 ( .A(n880), .B(n956), .CI(n896), .CO(n595), .S(n596) );
  CND2XL U2046 ( .A(n2063), .B(n2056), .Z(n1868) );
  CND2XL U2047 ( .A(n2063), .B(n2080), .Z(n1869) );
  CND2X1 U2048 ( .A(n2056), .B(n2080), .Z(n1870) );
  CND3X1 U2049 ( .A(n1868), .B(n1869), .C(n1870), .Z(n455) );
  CND2XL U2050 ( .A(n1581), .B(n1754), .Z(n1871) );
  CND2XL U2051 ( .A(n1754), .B(n455), .Z(n1873) );
  CND3X1 U2052 ( .A(n1871), .B(n1872), .C(n1873), .Z(n421) );
  CND2X2 U2053 ( .A(n1876), .B(n1877), .Z(n1944) );
  CIVXL U2054 ( .A(n693), .Z(n1874) );
  CND2XL U2055 ( .A(n529), .B(n2138), .Z(n1878) );
  CND2XL U2056 ( .A(n529), .B(n527), .Z(n1879) );
  CND2XL U2057 ( .A(n2138), .B(n527), .Z(n1880) );
  CND3X1 U2058 ( .A(n1878), .B(n1879), .C(n1880), .Z(n499) );
  CND3X2 U2059 ( .A(n2195), .B(n2196), .C(n2197), .Z(n539) );
  CIVX1 U2060 ( .A(n194), .Z(n192) );
  CEOX2 U2061 ( .A(n1071), .B(n941), .Z(n1881) );
  CEOX2 U2062 ( .A(n1806), .B(n1881), .Z(n712) );
  CND3X1 U2063 ( .A(n1882), .B(n1883), .C(n1884), .Z(n711) );
  CEOXL U2064 ( .A(n1885), .B(n532), .Z(n522) );
  CND2XL U2065 ( .A(n532), .B(n551), .Z(n1886) );
  CND2XL U2066 ( .A(n532), .B(n549), .Z(n1887) );
  CND3XL U2067 ( .A(n1886), .B(n1887), .C(n1888), .Z(n521) );
  CEOX1 U2068 ( .A(n931), .B(n877), .Z(n1889) );
  CND2XL U2069 ( .A(n863), .B(n877), .Z(n1890) );
  CND2XL U2070 ( .A(n863), .B(n931), .Z(n1891) );
  CND2XL U2071 ( .A(n877), .B(n931), .Z(n1892) );
  CND3XL U2072 ( .A(n1890), .B(n1891), .C(n1892), .Z(n531) );
  CFA1XL U2073 ( .A(n878), .B(n954), .CI(n912), .CO(n551), .S(n552) );
  CENXL U2074 ( .A(n1388), .B(n2002), .Z(n1166) );
  CENXL U2075 ( .A(n2208), .B(n1698), .Z(n1172) );
  CENXL U2076 ( .A(n1389), .B(n1698), .Z(n1167) );
  CENXL U2077 ( .A(n1396), .B(n1698), .Z(n1174) );
  CENXL U2078 ( .A(n2203), .B(n1560), .Z(n1178) );
  CEOX4 U2079 ( .A(n2234), .B(a[6]), .Z(n2029) );
  CENXL U2080 ( .A(n2234), .B(n2207), .Z(n1298) );
  CENXL U2081 ( .A(n2234), .B(n1396), .Z(n1299) );
  CND2X2 U2082 ( .A(net179371), .B(n1985), .Z(n1987) );
  CIVX8 U2083 ( .A(n2032), .Z(n42) );
  CEO3X2 U2084 ( .A(n2050), .B(n2045), .C(n2071), .Z(n528) );
  CND2X1 U2085 ( .A(n2050), .B(n2045), .Z(n1893) );
  CND2X1 U2086 ( .A(n2050), .B(n2071), .Z(n1894) );
  CND2X1 U2087 ( .A(n2045), .B(n2071), .Z(n1895) );
  CND3X2 U2088 ( .A(n1893), .B(n1894), .C(n1895), .Z(n527) );
  CND2XL U2089 ( .A(n1696), .B(n2139), .Z(n1896) );
  CND2X1 U2090 ( .A(n2139), .B(n528), .Z(n1898) );
  CEOX1 U2091 ( .A(n1041), .B(n987), .Z(n1899) );
  CND2XL U2092 ( .A(n1697), .B(n987), .Z(n1900) );
  CND2XL U2093 ( .A(n1697), .B(n1041), .Z(n1901) );
  CND2XL U2094 ( .A(n987), .B(n1041), .Z(n1902) );
  CND3X1 U2095 ( .A(n1900), .B(n1901), .C(n1902), .Z(n709) );
  COND2XL U2096 ( .A(n18), .B(n1327), .C(n1326), .D(n2185), .Z(n1041) );
  CIVXL U2097 ( .A(n208), .Z(n1903) );
  COND2X1 U2098 ( .A(n53), .B(n1223), .C(n50), .D(n1222), .Z(n941) );
  CENX1 U2099 ( .A(n2202), .B(n1975), .Z(n1223) );
  COND2XL U2100 ( .A(n2190), .B(n1138), .C(n1693), .D(n1137), .Z(n860) );
  COND2XL U2101 ( .A(n1904), .B(n1135), .C(n1864), .D(n1134), .Z(n857) );
  COND2XL U2102 ( .A(n2190), .B(n1144), .C(n1693), .D(n1143), .Z(n866) );
  COND2XL U2103 ( .A(n1904), .B(n1137), .C(n1693), .D(n1136), .Z(n859) );
  COND2XL U2104 ( .A(n2190), .B(n1136), .C(n1864), .D(n1135), .Z(n858) );
  CENXL U2105 ( .A(n1975), .B(n1385), .Z(n1207) );
  CENXL U2106 ( .A(n2205), .B(n1975), .Z(n1220) );
  CENXL U2107 ( .A(n2204), .B(n1975), .Z(n1221) );
  CENXL U2108 ( .A(net33480), .B(n2255), .Z(n1202) );
  COR2X2 U2109 ( .A(n536), .B(n557), .Z(n2015) );
  CENX1 U2110 ( .A(n573), .B(n2130), .Z(n2027) );
  CND3X2 U2111 ( .A(n1981), .B(n1982), .C(n1983), .Z(n573) );
  CND2XL U2112 ( .A(n1412), .B(n1864), .Z(n1904) );
  CEO3X2 U2113 ( .A(n710), .B(n708), .C(n719), .Z(n704) );
  CEOX2 U2114 ( .A(n706), .B(n717), .Z(n1906) );
  CEOX2 U2115 ( .A(n1906), .B(n704), .Z(n702) );
  CND2X1 U2116 ( .A(n710), .B(n708), .Z(n1907) );
  CND2X1 U2117 ( .A(n710), .B(n719), .Z(n1908) );
  CND2X1 U2118 ( .A(n708), .B(n719), .Z(n1909) );
  CND3X2 U2119 ( .A(n1907), .B(n1908), .C(n1909), .Z(n703) );
  CND2XL U2120 ( .A(n706), .B(n717), .Z(n1910) );
  CND2XL U2121 ( .A(n706), .B(n704), .Z(n1911) );
  CND2XL U2122 ( .A(n717), .B(n704), .Z(n1912) );
  CND3XL U2123 ( .A(n1910), .B(n1911), .C(n1912), .Z(n701) );
  CEOX1 U2124 ( .A(n695), .B(n697), .Z(n1913) );
  CND2X1 U2125 ( .A(n699), .B(n697), .Z(n1914) );
  CND2X1 U2126 ( .A(n699), .B(n695), .Z(n1915) );
  CND2X1 U2127 ( .A(n697), .B(n695), .Z(n1916) );
  CND3X1 U2128 ( .A(n1914), .B(n1915), .C(n1916), .Z(n677) );
  CNIVX2 U2129 ( .A(n700), .Z(n1917) );
  CND2X1 U2130 ( .A(n467), .B(n469), .Z(net180105) );
  CND2X1 U2131 ( .A(n467), .B(n446), .Z(net180106) );
  COND2XL U2132 ( .A(n44), .B(n1236), .C(n1235), .D(n42), .Z(n953) );
  CND2XL U2133 ( .A(n700), .B(n696), .Z(n1928) );
  CIVXL U2134 ( .A(n468), .Z(net180094) );
  CFA1XL U2135 ( .A(n898), .B(n1036), .CI(n916), .CO(n633), .S(n634) );
  CND2XL U2136 ( .A(n545), .B(n524), .Z(n1921) );
  CND2XL U2137 ( .A(n545), .B(n2137), .Z(n1922) );
  CND2XL U2138 ( .A(n524), .B(n2137), .Z(n1923) );
  CND3XL U2139 ( .A(n1921), .B(n1922), .C(n1923), .Z(n517) );
  CND2X1 U2140 ( .A(n2192), .B(n2191), .Z(n1924) );
  CND2X2 U2141 ( .A(n2193), .B(n1925), .Z(n545) );
  CIVX2 U2142 ( .A(n1924), .Z(n1925) );
  CND2XL U2143 ( .A(n2127), .B(n2130), .Z(n2191) );
  CND3XL U2144 ( .A(net180016), .B(net180017), .C(net180018), .Z(n419) );
  CENXL U2145 ( .A(net33480), .B(n2002), .Z(n1181) );
  CEOX2 U2146 ( .A(n696), .B(n698), .Z(n1926) );
  CEOX2 U2147 ( .A(n1926), .B(n1917), .Z(n692) );
  CND2XL U2148 ( .A(n700), .B(n698), .Z(n1927) );
  CND2XL U2149 ( .A(n698), .B(n696), .Z(n1929) );
  CND3X1 U2150 ( .A(n1927), .B(n1928), .C(n1929), .Z(n691) );
  CND3X1 U2151 ( .A(n1930), .B(n1931), .C(n1932), .Z(n459) );
  CNR2XL U2152 ( .A(net179834), .B(n487), .Z(n1938) );
  CEO3X1 U2153 ( .A(n466), .B(n1960), .C(n489), .Z(net179834) );
  COND2XL U2154 ( .A(n2190), .B(n1142), .C(n1693), .D(n1141), .Z(n864) );
  COND2XL U2155 ( .A(n2190), .B(n1140), .C(n1864), .D(n1139), .Z(n862) );
  CENX1 U2156 ( .A(n1396), .B(n2216), .Z(n1123) );
  CIVX1 U2157 ( .A(n186), .Z(n185) );
  CIVXL U2158 ( .A(n1597), .Z(n338) );
  CND3X1 U2159 ( .A(n1945), .B(n1946), .C(n1947), .Z(n675) );
  CNR2X2 U2160 ( .A(n1939), .B(n188), .Z(n186) );
  COND1X1 U2161 ( .A(n206), .B(n189), .C(n190), .Z(n188) );
  CND2X2 U2162 ( .A(n2020), .B(n2015), .Z(n189) );
  CIVXL U2163 ( .A(net180475), .Z(net179912) );
  CIVXL U2164 ( .A(net179912), .Z(net179913) );
  CND2X1 U2165 ( .A(n1985), .B(n1778), .Z(n1942) );
  CND2XL U2166 ( .A(n104), .B(n1940), .Z(n1943) );
  CIVXL U2167 ( .A(n1814), .Z(n1941) );
  CND2X2 U2168 ( .A(n1408), .B(n105), .Z(n107) );
  CND2XL U2169 ( .A(n682), .B(n1614), .Z(n1945) );
  CND2XL U2170 ( .A(n693), .B(n684), .Z(n1947) );
  COR2X1 U2171 ( .A(n1164), .B(n1970), .Z(n1948) );
  COR2X1 U2172 ( .A(n74), .B(n1163), .Z(n1949) );
  CND2X2 U2173 ( .A(n1948), .B(n1949), .Z(n885) );
  CENX1 U2174 ( .A(net33082), .B(n1969), .Z(n1164) );
  CND2XL U2175 ( .A(n816), .B(n1674), .Z(n1950) );
  CND2XL U2176 ( .A(n1674), .B(n846), .Z(n1952) );
  CND3XL U2177 ( .A(n1950), .B(n1951), .C(n1952), .Z(n405) );
  COND2X1 U2178 ( .A(n1964), .B(n1123), .C(n89), .D(n1122), .Z(n846) );
  CEOX1 U2179 ( .A(n2142), .B(n523), .Z(n1953) );
  CND2X1 U2180 ( .A(n500), .B(n523), .Z(n1954) );
  CND2X1 U2181 ( .A(n523), .B(n2142), .Z(n1956) );
  CND3X2 U2182 ( .A(n1954), .B(n1955), .C(n1956), .Z(n493) );
  CND2X1 U2183 ( .A(n2067), .B(n2078), .Z(n1957) );
  CIVXL U2184 ( .A(n1938), .Z(n337) );
  CNR2IX1 U2185 ( .B(net33082), .A(n1652), .Z(n924) );
  COND2X1 U2186 ( .A(n36), .B(n1276), .C(n1275), .D(n33), .Z(n992) );
  COND2X1 U2187 ( .A(n36), .B(n1274), .C(n1273), .D(n33), .Z(n990) );
  COND2X1 U2188 ( .A(n36), .B(n1270), .C(n1269), .D(n33), .Z(n986) );
  COND2X1 U2189 ( .A(n36), .B(n1272), .C(n1271), .D(n33), .Z(n988) );
  CENXL U2190 ( .A(n2205), .B(n1694), .Z(n1140) );
  CIVX1 U2191 ( .A(n2244), .Z(n2239) );
  CIVX4 U2192 ( .A(n30), .Z(n2244) );
  CENXL U2193 ( .A(n2232), .B(n2202), .Z(n1304) );
  CENXL U2194 ( .A(n2232), .B(n2204), .Z(n1302) );
  CENXL U2195 ( .A(n2232), .B(n2203), .Z(n1303) );
  CENXL U2196 ( .A(n2232), .B(n2205), .Z(n1301) );
  CFA1X1 U2197 ( .A(n932), .B(n842), .CI(n894), .CO(n553), .S(n554) );
  CND2X2 U2198 ( .A(n1409), .B(n1984), .Z(n102) );
  CND2X1 U2199 ( .A(n1995), .B(n1996), .Z(n1409) );
  CENXL U2200 ( .A(n2203), .B(n1752), .Z(n1142) );
  CENX4 U2201 ( .A(n2247), .B(a[10]), .Z(n50) );
  CENXL U2202 ( .A(n2238), .B(b[25]), .Z(n1254) );
  CENXL U2203 ( .A(n2241), .B(n2206), .Z(n1271) );
  CENXL U2204 ( .A(n2242), .B(net33482), .Z(n1278) );
  CFA1X1 U2205 ( .A(n1073), .B(n943), .CI(n1015), .CO(n735), .S(n736) );
  CENXL U2206 ( .A(n2227), .B(n2206), .Z(n1331) );
  CENXL U2207 ( .A(n2227), .B(n1396), .Z(n1330) );
  CENXL U2208 ( .A(n2227), .B(n2207), .Z(n1329) );
  CENXL U2209 ( .A(n2227), .B(n1387), .Z(n1321) );
  CFA1X1 U2210 ( .A(n967), .B(n1075), .CI(n1045), .CO(n755), .S(n756) );
  COND2X1 U2211 ( .A(n18), .B(n1331), .C(n1330), .D(n2185), .Z(n1045) );
  CENXL U2212 ( .A(n142), .B(n1627), .Z(product[8]) );
  COND2XL U2213 ( .A(n27), .B(n1288), .C(n1287), .D(n2009), .Z(n1003) );
  COND2XL U2214 ( .A(n27), .B(n1291), .C(n1290), .D(n2009), .Z(n1006) );
  COND2XL U2215 ( .A(n27), .B(n1287), .C(n1286), .D(n2009), .Z(n1002) );
  COND2XL U2216 ( .A(n27), .B(n1285), .C(n1284), .D(n2009), .Z(n1000) );
  COND2XL U2217 ( .A(n27), .B(n1294), .C(n1293), .D(n2009), .Z(n1009) );
  COND2XL U2218 ( .A(n27), .B(n1293), .C(n1292), .D(n2009), .Z(n1008) );
  COND2XL U2219 ( .A(n27), .B(n1295), .C(n1294), .D(n2009), .Z(n1010) );
  COND2XL U2220 ( .A(n27), .B(n1299), .C(n1298), .D(n2009), .Z(n1014) );
  COND2XL U2221 ( .A(n27), .B(n1297), .C(n1296), .D(n2009), .Z(n1012) );
  COND2X1 U2222 ( .A(n1964), .B(n1128), .C(n1127), .D(n89), .Z(n851) );
  COND2X1 U2223 ( .A(n1964), .B(n1692), .C(n89), .D(n1128), .Z(n852) );
  CND2X2 U2224 ( .A(n1979), .B(n1980), .Z(n1412) );
  CND2X2 U2225 ( .A(a[18]), .B(n1978), .Z(n1979) );
  CIVXL U2226 ( .A(n1669), .Z(n1961) );
  CIVXL U2227 ( .A(n1961), .Z(n1962) );
  COND2X1 U2228 ( .A(n18), .B(n1336), .C(n1335), .D(n2185), .Z(n1050) );
  CNR2X2 U2229 ( .A(n189), .B(n205), .Z(n187) );
  CND2X2 U2230 ( .A(n2017), .B(n342), .Z(n205) );
  CND2IXL U2231 ( .B(net33082), .A(n2218), .Z(n1109) );
  CENXL U2232 ( .A(net33080), .B(n2218), .Z(n1108) );
  CENXL U2233 ( .A(n2205), .B(n2218), .Z(n1101) );
  CENXL U2234 ( .A(n2203), .B(n2218), .Z(n1103) );
  CENXL U2235 ( .A(n2202), .B(n2218), .Z(n1104) );
  CENXL U2236 ( .A(n2201), .B(n2218), .Z(n1105) );
  CENXL U2237 ( .A(net33480), .B(n2218), .Z(n1106) );
  CENXL U2238 ( .A(net33482), .B(n2218), .Z(n1107) );
  CENXL U2239 ( .A(n2204), .B(n2218), .Z(n1102) );
  CNIVX3 U2240 ( .A(n99), .Z(n2218) );
  CIVXL U2241 ( .A(net179544), .Z(net179686) );
  CIVXL U2242 ( .A(n1621), .Z(n1435) );
  CENXL U2243 ( .A(net179680), .B(n164), .Z(product[29]) );
  CNR2IX1 U2244 ( .B(net33082), .A(n50), .Z(n946) );
  CANR1X1 U2245 ( .A(n232), .B(n2021), .C(n227), .Z(n225) );
  COND2XL U2246 ( .A(n36), .B(n1257), .C(n1256), .D(n33), .Z(n973) );
  COND2XL U2247 ( .A(n36), .B(n1263), .C(n1262), .D(n33), .Z(n979) );
  COND2XL U2248 ( .A(n36), .B(n1255), .C(n1254), .D(n33), .Z(n971) );
  COND2XL U2249 ( .A(n36), .B(n1265), .C(n1264), .D(n33), .Z(n981) );
  COND2XL U2250 ( .A(n36), .B(n1266), .C(n1265), .D(n33), .Z(n982) );
  COND2XL U2251 ( .A(n36), .B(n1256), .C(n1255), .D(n33), .Z(n972) );
  COND2XL U2252 ( .A(n36), .B(n1258), .C(n1257), .D(n33), .Z(n974) );
  COND2XL U2253 ( .A(n36), .B(n1264), .C(n1263), .D(n33), .Z(n980) );
  COND2XL U2254 ( .A(n36), .B(n1261), .C(n1260), .D(n33), .Z(n977) );
  COND2XL U2255 ( .A(n36), .B(n1260), .C(n1259), .D(n33), .Z(n976) );
  COND2XL U2256 ( .A(n36), .B(n1259), .C(n1258), .D(n33), .Z(n975) );
  COND2XL U2257 ( .A(n36), .B(n1262), .C(n1261), .D(n33), .Z(n978) );
  COND2XL U2258 ( .A(n36), .B(n1268), .C(n1267), .D(n33), .Z(n984) );
  COND2XL U2259 ( .A(n36), .B(n1267), .C(n1266), .D(n33), .Z(n983) );
  COND2XL U2260 ( .A(n36), .B(n1269), .C(n1268), .D(n33), .Z(n985) );
  COND2XL U2261 ( .A(n36), .B(n1275), .C(n1274), .D(n33), .Z(n991) );
  COND2XL U2262 ( .A(n1279), .B(n36), .C(n1278), .D(n33), .Z(n995) );
  COND2XL U2263 ( .A(n36), .B(n1271), .C(n1270), .D(n33), .Z(n987) );
  COND2XL U2264 ( .A(n36), .B(n2243), .C(n33), .D(n1280), .Z(n811) );
  COR2XL U2265 ( .A(n1436), .B(n1964), .Z(n1977) );
  CANR1X1 U2266 ( .A(n201), .B(n1936), .C(n192), .Z(n190) );
  CANR1X1 U2267 ( .A(n338), .B(n185), .C(n182), .Z(n180) );
  CANR1XL U2268 ( .A(n297), .B(n2014), .C(n292), .Z(n290) );
  CND2X1 U2269 ( .A(n1988), .B(n1989), .Z(n100) );
  COND2X1 U2270 ( .A(n9), .B(n1369), .C(n6), .D(n1368), .Z(n1082) );
  COND1X1 U2271 ( .A(n317), .B(n315), .C(n316), .Z(n314) );
  CNR2XL U2272 ( .A(n792), .B(n795), .Z(n315) );
  CANR1X1 U2273 ( .A(n322), .B(n2023), .C(n319), .Z(n317) );
  CND2IXL U2274 ( .B(net33082), .A(n1621), .Z(n1120) );
  CENXL U2275 ( .A(n2204), .B(n2217), .Z(n1113) );
  CENXL U2276 ( .A(n2203), .B(n2217), .Z(n1114) );
  CENXL U2277 ( .A(n2202), .B(n2217), .Z(n1115) );
  CENXL U2278 ( .A(n2201), .B(n1621), .Z(n1116) );
  CENXL U2279 ( .A(n1396), .B(n2217), .Z(n1110) );
  CENXL U2280 ( .A(net33080), .B(n2217), .Z(n1119) );
  CND2X2 U2281 ( .A(n1407), .B(n110), .Z(n112) );
  CND2IX1 U2282 ( .B(n2006), .A(n74), .Z(n1970) );
  CFA1X1 U2283 ( .A(n904), .B(n922), .CI(n942), .CO(n725), .S(n726) );
  COND2X1 U2284 ( .A(n18), .B(n1333), .C(n1332), .D(n2185), .Z(n1047) );
  CIVXL U2285 ( .A(n1652), .Z(n1967) );
  CIVX2 U2286 ( .A(n1967), .Z(n1968) );
  COND2XL U2287 ( .A(n9), .B(n1348), .C(n6), .D(n1347), .Z(n1061) );
  CND2IXL U2288 ( .B(net33082), .A(n1814), .Z(n1100) );
  CENXL U2289 ( .A(net33080), .B(n1814), .Z(n1099) );
  CENXL U2290 ( .A(n2203), .B(n1814), .Z(n1094) );
  CENXL U2291 ( .A(net33480), .B(n104), .Z(n1097) );
  CENXL U2292 ( .A(n2202), .B(n104), .Z(n1095) );
  CENXL U2293 ( .A(n2201), .B(n104), .Z(n1096) );
  CENXL U2294 ( .A(net33482), .B(n104), .Z(n1098) );
  CNIVX4 U2295 ( .A(n71), .Z(n1969) );
  COND2X1 U2296 ( .A(n1226), .B(n53), .C(n1225), .D(n50), .Z(n944) );
  COND2XL U2297 ( .A(n2190), .B(n1139), .C(n1864), .D(n1138), .Z(n861) );
  CENXL U2298 ( .A(n2208), .B(n1606), .Z(n1121) );
  CENXL U2299 ( .A(n2204), .B(n1606), .Z(n1126) );
  CENXL U2300 ( .A(n2205), .B(n1755), .Z(n1125) );
  CENXL U2301 ( .A(n2207), .B(n1755), .Z(n1122) );
  CENXL U2302 ( .A(net33080), .B(n1755), .Z(n1132) );
  CENXL U2303 ( .A(n1755), .B(net33482), .Z(n1131) );
  CENXL U2304 ( .A(n2202), .B(n1755), .Z(n1128) );
  CENXL U2305 ( .A(n2203), .B(n1755), .Z(n1127) );
  CENXL U2306 ( .A(net33480), .B(n1755), .Z(n1130) );
  CENXL U2307 ( .A(n2210), .B(n1694), .Z(n1134) );
  CENXL U2308 ( .A(n1396), .B(n1752), .Z(n1138) );
  CENXL U2309 ( .A(n2207), .B(n1752), .Z(n1137) );
  CENXL U2310 ( .A(n2209), .B(n1752), .Z(n1135) );
  CENXL U2311 ( .A(n2206), .B(n1752), .Z(n1139) );
  CENXL U2312 ( .A(n2208), .B(n1752), .Z(n1136) );
  CENXL U2313 ( .A(n2202), .B(n2215), .Z(n1143) );
  CENXL U2314 ( .A(net33080), .B(n2215), .Z(n1147) );
  CENXL U2315 ( .A(n2204), .B(n1752), .Z(n1141) );
  COND2X1 U2316 ( .A(n53), .B(n1224), .C(n1223), .D(n50), .Z(n942) );
  CIVXL U2317 ( .A(n1969), .Z(n1438) );
  COND2XL U2318 ( .A(n107), .B(n1096), .C(n105), .D(n1095), .Z(n822) );
  COND2XL U2319 ( .A(n107), .B(n1097), .C(n105), .D(n1096), .Z(n823) );
  COND2XL U2320 ( .A(n1099), .B(n107), .C(n105), .D(n1098), .Z(n825) );
  COND2X1 U2321 ( .A(n1805), .B(n1100), .C(n1941), .D(n107), .Z(n801) );
  COND2X1 U2322 ( .A(n1807), .B(n1093), .C(net179686), .D(n112), .Z(n800) );
  COND2XL U2323 ( .A(n77), .B(n1153), .C(n74), .D(n1152), .Z(n874) );
  COND2XL U2324 ( .A(n77), .B(n1151), .C(n74), .D(n1150), .Z(n872) );
  COND2XL U2325 ( .A(n77), .B(n1150), .C(n74), .D(n1149), .Z(n871) );
  COND2XL U2326 ( .A(n77), .B(n1154), .C(n74), .D(n1153), .Z(n875) );
  COND2XL U2327 ( .A(n77), .B(n1155), .C(n74), .D(n1154), .Z(n876) );
  COND2XL U2328 ( .A(n77), .B(n1160), .C(n74), .D(n1159), .Z(n881) );
  COND2XL U2329 ( .A(n77), .B(n1159), .C(n74), .D(n1158), .Z(n880) );
  COND2XL U2330 ( .A(n77), .B(n1152), .C(n74), .D(n1151), .Z(n873) );
  CENXL U2331 ( .A(n2201), .B(net179544), .Z(n1089) );
  CENXL U2332 ( .A(net33080), .B(net179544), .Z(n1092) );
  COND2XL U2333 ( .A(n1619), .B(n1194), .C(n1193), .D(n1968), .Z(n913) );
  COND2XL U2334 ( .A(n1619), .B(n1188), .C(n1187), .D(n1968), .Z(n907) );
  COND2XL U2335 ( .A(n1619), .B(n1191), .C(n1190), .D(n1968), .Z(n910) );
  COND2XL U2336 ( .A(n1619), .B(n1192), .C(n1191), .D(n1968), .Z(n911) );
  COND2XL U2337 ( .A(n1619), .B(n1189), .C(n1188), .D(n1968), .Z(n908) );
  COND2XL U2338 ( .A(n1619), .B(n1190), .C(n1189), .D(n1968), .Z(n909) );
  COND2XL U2339 ( .A(n1619), .B(n1187), .C(n1186), .D(n1968), .Z(n906) );
  COND2XL U2340 ( .A(n1619), .B(n1186), .C(n1185), .D(n1968), .Z(n905) );
  COND2XL U2341 ( .A(n1619), .B(n1196), .C(n1195), .D(n1968), .Z(n915) );
  COND2XL U2342 ( .A(n1619), .B(n1195), .C(n1194), .D(n1968), .Z(n914) );
  COND2XL U2343 ( .A(n1619), .B(n1198), .C(n1968), .D(n1197), .Z(n917) );
  COND2XL U2344 ( .A(n1619), .B(n1193), .C(n1192), .D(n1652), .Z(n912) );
  COND2XL U2345 ( .A(n1619), .B(n1197), .C(n1196), .D(n1652), .Z(n916) );
  COND2XL U2346 ( .A(n61), .B(n1199), .C(n1652), .D(n1198), .Z(n918) );
  COND2XL U2347 ( .A(n61), .B(n1200), .C(n1652), .D(n1199), .Z(n919) );
  COND2XL U2348 ( .A(n61), .B(n1201), .C(n1652), .D(n1200), .Z(n920) );
  COND2XL U2349 ( .A(n1204), .B(n61), .C(n1652), .D(n1203), .Z(n923) );
  COND2XL U2350 ( .A(n1623), .B(n1172), .C(n1607), .D(n1171), .Z(n892) );
  COND2XL U2351 ( .A(n1623), .B(n1173), .C(n1607), .D(n1172), .Z(n893) );
  COND2XL U2352 ( .A(n69), .B(n1180), .C(n1607), .D(n1179), .Z(n900) );
  COND2X1 U2353 ( .A(n69), .B(n1561), .C(n66), .D(n1184), .Z(n807) );
  COND2XL U2354 ( .A(n1676), .B(n1127), .C(n1617), .D(n1126), .Z(n850) );
  COND2XL U2355 ( .A(n69), .B(n1178), .C(n1607), .D(n1177), .Z(n898) );
  COND2XL U2356 ( .A(n1623), .B(n1179), .C(n1607), .D(n1178), .Z(n899) );
  CNR2X1 U2357 ( .A(n183), .B(n1937), .Z(n172) );
  CENX2 U2358 ( .A(a[16]), .B(n2214), .Z(n2006) );
  COND2XL U2359 ( .A(n77), .B(n1156), .C(n74), .D(n1155), .Z(n877) );
  COND2XL U2360 ( .A(n77), .B(n1157), .C(n74), .D(n1156), .Z(n878) );
  COND2XL U2361 ( .A(n77), .B(n1158), .C(n74), .D(n1157), .Z(n879) );
  COND2XL U2362 ( .A(n77), .B(n1162), .C(n74), .D(n1161), .Z(n883) );
  COND2XL U2363 ( .A(n1676), .B(n1125), .C(n1617), .D(n1124), .Z(n848) );
  CIVX4 U2364 ( .A(n2222), .Z(n2220) );
  CIVX3 U2365 ( .A(n3), .Z(n2222) );
  CENXL U2366 ( .A(n120), .B(n157), .Z(product[30]) );
  CNR2IX1 U2367 ( .B(net33082), .A(n74), .Z(n886) );
  CENXL U2368 ( .A(n2212), .B(n1969), .Z(n1149) );
  CENXL U2369 ( .A(n2211), .B(n1969), .Z(n1150) );
  CENXL U2370 ( .A(n2208), .B(n1969), .Z(n1153) );
  CENXL U2371 ( .A(n2207), .B(n1969), .Z(n1154) );
  CENXL U2372 ( .A(n2203), .B(n1969), .Z(n1159) );
  CENXL U2373 ( .A(n2209), .B(n1969), .Z(n1152) );
  CENXL U2374 ( .A(n2210), .B(n1969), .Z(n1151) );
  CENXL U2375 ( .A(n2204), .B(n1969), .Z(n1158) );
  CENXL U2376 ( .A(n2205), .B(n1969), .Z(n1157) );
  CENXL U2377 ( .A(n2201), .B(n1969), .Z(n1161) );
  CENXL U2378 ( .A(n1396), .B(n1969), .Z(n1155) );
  CENXL U2379 ( .A(n2206), .B(n1969), .Z(n1156) );
  CENXL U2380 ( .A(n2202), .B(n1969), .Z(n1160) );
  CENX4 U2381 ( .A(n1752), .B(a[20]), .Z(n89) );
  CND2X2 U2382 ( .A(n1972), .B(n1833), .Z(n1974) );
  CND2X2 U2383 ( .A(n1973), .B(n1974), .Z(n95) );
  CIVXL U2384 ( .A(n1755), .Z(n1972) );
  COND2XL U2385 ( .A(n1111), .B(n1669), .C(n95), .D(n1110), .Z(n835) );
  COND2XL U2386 ( .A(n1962), .B(n1116), .C(n95), .D(n1115), .Z(n840) );
  COND2XL U2387 ( .A(n1962), .B(n1114), .C(n95), .D(n1113), .Z(n838) );
  COND2XL U2388 ( .A(n1669), .B(n1115), .C(n95), .D(n1114), .Z(n839) );
  COND2XL U2389 ( .A(n1669), .B(n1113), .C(n95), .D(n1112), .Z(n837) );
  CNIVX4 U2390 ( .A(n48), .Z(n1975) );
  COR2XL U2391 ( .A(n1133), .B(n89), .Z(n1976) );
  CND2IXL U2392 ( .B(net33082), .A(n1755), .Z(n1133) );
  CIVXL U2393 ( .A(n2216), .Z(n1436) );
  CND2X1 U2394 ( .A(n2052), .B(n2049), .Z(n1981) );
  CND2X1 U2395 ( .A(n2052), .B(n2070), .Z(n1982) );
  CND2X1 U2396 ( .A(n2049), .B(n2070), .Z(n1983) );
  CND2XL U2397 ( .A(n2130), .B(n573), .Z(n2193) );
  CND2XL U2398 ( .A(n2127), .B(n573), .Z(n2192) );
  COND1X1 U2399 ( .A(n241), .B(n224), .C(n225), .Z(n223) );
  CENXL U2400 ( .A(n2209), .B(n1698), .Z(n1171) );
  CENXL U2401 ( .A(n2210), .B(n1698), .Z(n1170) );
  CENXL U2402 ( .A(n2212), .B(n1698), .Z(n1168) );
  CENXL U2403 ( .A(n2205), .B(n1560), .Z(n1176) );
  CENXL U2404 ( .A(n2202), .B(n2002), .Z(n1179) );
  CENXL U2405 ( .A(n2254), .B(n1387), .Z(n1186) );
  CENXL U2406 ( .A(n2254), .B(n1388), .Z(n1187) );
  CENXL U2407 ( .A(n2254), .B(n1389), .Z(n1188) );
  CENXL U2408 ( .A(n2254), .B(n1386), .Z(n1185) );
  CENXL U2409 ( .A(n2254), .B(n2212), .Z(n1189) );
  CENXL U2410 ( .A(n2254), .B(n2211), .Z(n1190) );
  CENXL U2411 ( .A(n2210), .B(n2254), .Z(n1191) );
  CENXL U2412 ( .A(n2204), .B(n2254), .Z(n1198) );
  CENXL U2413 ( .A(n2203), .B(n2254), .Z(n1199) );
  CENXL U2414 ( .A(n2202), .B(n2254), .Z(n1200) );
  CENXL U2415 ( .A(n2201), .B(n2254), .Z(n1201) );
  CND2X2 U2416 ( .A(n1986), .B(n1987), .Z(n110) );
  COND2XL U2417 ( .A(n112), .B(n1091), .C(n1090), .D(n1807), .Z(n818) );
  COND2XL U2418 ( .A(n112), .B(n1092), .C(n110), .D(n1091), .Z(n819) );
  COND2XL U2419 ( .A(n112), .B(n1090), .C(n110), .D(n1089), .Z(n817) );
  COND2XL U2420 ( .A(n1120), .B(n95), .C(n1435), .D(n1669), .Z(n803) );
  CND2XL U2421 ( .A(a[24]), .B(n2217), .Z(n1988) );
  CIVXL U2422 ( .A(n167), .Z(n336) );
  COND2XL U2423 ( .A(n1117), .B(n1962), .C(n95), .D(n1116), .Z(n841) );
  CIVXL U2424 ( .A(n162), .Z(n335) );
  CNIVX4 U2425 ( .A(n86), .Z(n2216) );
  CND2XL U2426 ( .A(a[24]), .B(n1994), .Z(n1995) );
  CND2XL U2427 ( .A(n1993), .B(n2218), .Z(n1996) );
  COND2XL U2428 ( .A(n1108), .B(n102), .C(n1984), .D(n1107), .Z(n833) );
  COND2XL U2429 ( .A(n1106), .B(n102), .C(n1984), .D(n1105), .Z(n831) );
  COND2XL U2430 ( .A(n1105), .B(n102), .C(n1984), .D(n1104), .Z(n830) );
  COND2XL U2431 ( .A(n1104), .B(n102), .C(n1984), .D(n1103), .Z(n829) );
  COND2XL U2432 ( .A(n1103), .B(n102), .C(n1984), .D(n1102), .Z(n828) );
  COND2XL U2433 ( .A(n102), .B(n1102), .C(n1984), .D(n1101), .Z(n827) );
  CNIVX3 U2434 ( .A(n1399), .Z(n2204) );
  COR2XL U2435 ( .A(n1084), .B(n1054), .Z(n2024) );
  CNR2IXL U2436 ( .B(net33082), .A(n2009), .Z(n1024) );
  CENX1 U2437 ( .A(n2233), .B(net33480), .Z(n1306) );
  CENX1 U2438 ( .A(n2233), .B(net33482), .Z(n1307) );
  COAN1X1 U2439 ( .A(n301), .B(n289), .C(n1966), .Z(n2003) );
  COR2XL U2440 ( .A(n1306), .B(n2009), .Z(n2005) );
  COND1XL U2441 ( .A(n301), .B(n289), .C(n290), .Z(n288) );
  CND2X1 U2442 ( .A(n760), .B(n767), .Z(n294) );
  CIVX2 U2443 ( .A(n2250), .Z(n2247) );
  CNR2IXL U2444 ( .B(net33082), .A(n33), .Z(n996) );
  CENX2 U2445 ( .A(n12), .B(a[4]), .Z(n2009) );
  CENX1 U2446 ( .A(a[4]), .B(n2234), .Z(n2008) );
  CNIVX2 U2447 ( .A(n1393), .Z(n2209) );
  CNIVX2 U2448 ( .A(n1392), .Z(n2210) );
  COND2X1 U2449 ( .A(n97), .B(n1118), .C(n95), .D(n1117), .Z(n842) );
  CNR2XL U2450 ( .A(n1815), .B(n285), .Z(n280) );
  CNR2XL U2451 ( .A(n688), .B(n701), .Z(n254) );
  CNR2XL U2452 ( .A(n716), .B(n727), .Z(n271) );
  CND2XL U2453 ( .A(n702), .B(n715), .Z(n267) );
  CEOXL U2454 ( .A(n123), .B(n180), .Z(product[27]) );
  CND2XL U2455 ( .A(n2016), .B(n299), .Z(n141) );
  CND2XL U2456 ( .A(n2018), .B(n305), .Z(n142) );
  CNR2IXL U2457 ( .B(n1662), .A(n167), .Z(n165) );
  CND2XL U2458 ( .A(n294), .B(n2014), .Z(n140) );
  CND2IXL U2459 ( .B(n1815), .A(n283), .Z(n138) );
  CND2XL U2460 ( .A(n2021), .B(n229), .Z(n129) );
  CANR1X1 U2461 ( .A(n219), .B(n1844), .C(n212), .Z(n206) );
  CIVX1 U2462 ( .A(n214), .Z(n212) );
  CND2IXL U2463 ( .B(n307), .A(n308), .Z(n143) );
  CND2IXL U2464 ( .B(n315), .A(n316), .Z(n145) );
  CND2XL U2465 ( .A(n2022), .B(n313), .Z(n144) );
  CND2XL U2466 ( .A(n2024), .B(n329), .Z(n148) );
  CND2XL U2467 ( .A(n2023), .B(n321), .Z(n146) );
  CND2XL U2468 ( .A(n207), .B(n2015), .Z(n196) );
  CND2XL U2469 ( .A(n740), .B(n749), .Z(n283) );
  CNR2XL U2470 ( .A(n728), .B(n739), .Z(n276) );
  CND2XL U2471 ( .A(n344), .B(n234), .Z(n130) );
  CEOX1 U2472 ( .A(n855), .B(n981), .Z(n2186) );
  CND2XL U2473 ( .A(n345), .B(n239), .Z(n131) );
  CND2XL U2474 ( .A(n798), .B(n1053), .Z(n324) );
  CND2XL U2475 ( .A(n792), .B(n795), .Z(n316) );
  COR2XL U2476 ( .A(n1085), .B(n814), .Z(n2007) );
  CND2IXL U2477 ( .B(net33082), .A(net179544), .Z(n1093) );
  COND2XL U2478 ( .A(n1623), .B(n1174), .C(n1607), .D(n1173), .Z(n894) );
  CIVX4 U2479 ( .A(n2033), .Z(n2185) );
  CEOXL U2480 ( .A(n835), .B(n871), .Z(n378) );
  CNIVX2 U2481 ( .A(n1390), .Z(n2212) );
  CNIVX2 U2482 ( .A(n1391), .Z(n2211) );
  CNIVX4 U2483 ( .A(n1401), .Z(n2202) );
  CNIVX4 U2484 ( .A(n1400), .Z(n2203) );
  CNIVX4 U2485 ( .A(n1398), .Z(n2205) );
  CNIVX4 U2486 ( .A(n1403), .Z(net33480) );
  CEO3X1 U2487 ( .A(n2010), .B(n2011), .C(n375), .Z(n370) );
  CEO3X1 U2488 ( .A(n2038), .B(n2088), .C(n2058), .Z(n2010) );
  CEO3X1 U2489 ( .A(n2077), .B(n2086), .C(n2036), .Z(n2011) );
  CEO3X1 U2490 ( .A(n2012), .B(n2166), .C(n395), .Z(n369) );
  CEO3X1 U2491 ( .A(n2051), .B(n2087), .C(n2047), .Z(n2012) );
  CENX1 U2492 ( .A(n204), .B(n126), .Z(product[24]) );
  CANR1XL U2493 ( .A(n2016), .B(n300), .C(n297), .Z(n295) );
  CENX1 U2494 ( .A(n141), .B(n300), .Z(product[9]) );
  CANR1XL U2495 ( .A(n280), .B(n288), .C(n281), .Z(n279) );
  COND1XL U2496 ( .A(n286), .B(n282), .C(n283), .Z(n281) );
  COND1XL U2497 ( .A(n285), .B(n2003), .C(n286), .Z(n284) );
  CANR1XL U2498 ( .A(n2015), .B(n208), .C(n201), .Z(n197) );
  CND2XL U2499 ( .A(n688), .B(n701), .Z(n255) );
  CND2XL U2500 ( .A(n716), .B(n727), .Z(n272) );
  COR2X1 U2501 ( .A(n715), .B(n702), .Z(n2013) );
  CANR1XL U2502 ( .A(n330), .B(n2024), .C(n327), .Z(n325) );
  CND2XL U2503 ( .A(n338), .B(n184), .Z(n124) );
  CENX1 U2504 ( .A(n215), .B(n127), .Z(product[23]) );
  COND1XL U2505 ( .A(n216), .B(n222), .C(n217), .Z(n215) );
  CENX1 U2506 ( .A(n144), .B(n314), .Z(product[6]) );
  CENX1 U2507 ( .A(n148), .B(n330), .Z(product[2]) );
  CENX1 U2508 ( .A(n146), .B(n322), .Z(product[4]) );
  CENX1 U2509 ( .A(n195), .B(n125), .Z(product[25]) );
  CND2XL U2510 ( .A(n1936), .B(n194), .Z(n125) );
  COND1XL U2511 ( .A(n196), .B(n222), .C(n197), .Z(n195) );
  CEOXL U2512 ( .A(n325), .B(n147), .Z(product[3]) );
  CND2X1 U2513 ( .A(n361), .B(n324), .Z(n147) );
  CEOXL U2514 ( .A(n128), .B(n222), .Z(product[22]) );
  CND2XL U2515 ( .A(n342), .B(n217), .Z(n128) );
  CEOX1 U2516 ( .A(n129), .B(n230), .Z(product[21]) );
  CANR1XL U2517 ( .A(n231), .B(n240), .C(n232), .Z(n230) );
  CND2X2 U2518 ( .A(n1410), .B(n95), .Z(n97) );
  COR2X1 U2519 ( .A(n767), .B(n760), .Z(n2014) );
  CND2X1 U2520 ( .A(n750), .B(n759), .Z(n286) );
  CND2X1 U2521 ( .A(n768), .B(n775), .Z(n299) );
  CND2X1 U2522 ( .A(n776), .B(n781), .Z(n305) );
  COR2X1 U2523 ( .A(n768), .B(n775), .Z(n2016) );
  COR2X1 U2524 ( .A(n558), .B(n579), .Z(n2017) );
  COR2X1 U2525 ( .A(n776), .B(n781), .Z(n2018) );
  CND2X1 U2526 ( .A(n558), .B(n579), .Z(n214) );
  CND2XL U2527 ( .A(n728), .B(n739), .Z(n277) );
  CEOX1 U2528 ( .A(n130), .B(n235), .Z(product[20]) );
  CANR1XL U2529 ( .A(n345), .B(n240), .C(n237), .Z(n235) );
  COND1XL U2530 ( .A(n239), .B(n233), .C(n234), .Z(n232) );
  CND2XL U2531 ( .A(n231), .B(n2021), .Z(n224) );
  CENX1 U2532 ( .A(n2019), .B(n538), .Z(n536) );
  CENX1 U2533 ( .A(n540), .B(n559), .Z(n2019) );
  COR2X1 U2534 ( .A(n535), .B(n512), .Z(n2020) );
  CNR2X1 U2535 ( .A(n488), .B(n511), .Z(n183) );
  CENX1 U2536 ( .A(n240), .B(n131), .Z(product[19]) );
  CNR2X1 U2537 ( .A(n782), .B(n787), .Z(n307) );
  CNR2X1 U2538 ( .A(n580), .B(n599), .Z(n216) );
  CNR2X1 U2539 ( .A(n798), .B(n1053), .Z(n323) );
  COR2X1 U2540 ( .A(n619), .B(n600), .Z(n2021) );
  CND2X1 U2541 ( .A(n580), .B(n599), .Z(n217) );
  CND3XL U2542 ( .A(n2187), .B(n2188), .C(n2189), .Z(n611) );
  CND2X1 U2543 ( .A(n1085), .B(n814), .Z(n332) );
  CND2X1 U2544 ( .A(n788), .B(n791), .Z(n313) );
  CND2X1 U2545 ( .A(n796), .B(n797), .Z(n321) );
  CND2X1 U2546 ( .A(n1084), .B(n1054), .Z(n329) );
  CND2X1 U2547 ( .A(n600), .B(n619), .Z(n229) );
  CND2X1 U2548 ( .A(n782), .B(n787), .Z(n308) );
  COR2X1 U2549 ( .A(n788), .B(n791), .Z(n2022) );
  COR2X1 U2550 ( .A(n796), .B(n797), .Z(n2023) );
  CENX1 U2551 ( .A(net33080), .B(n2229), .Z(n1339) );
  CNR2IX1 U2552 ( .B(net33082), .A(n42), .Z(n970) );
  CENX1 U2553 ( .A(n2225), .B(n2202), .Z(n1335) );
  CIVX2 U2554 ( .A(n2222), .Z(n2219) );
  CENX1 U2555 ( .A(n2239), .B(n2205), .Z(n1272) );
  CENX1 U2556 ( .A(n2236), .B(n2212), .Z(n1293) );
  CENX1 U2557 ( .A(n2248), .B(n2210), .Z(n1239) );
  CENX1 U2558 ( .A(n2248), .B(n2212), .Z(n1237) );
  CENX2 U2559 ( .A(n2254), .B(a[14]), .Z(n66) );
  CANR1XL U2560 ( .A(n261), .B(n242), .C(n243), .Z(n241) );
  CNR2X1 U2561 ( .A(n244), .B(n247), .Z(n242) );
  COND1XL U2562 ( .A(n244), .B(n248), .C(n245), .Z(n243) );
  CENX1 U2563 ( .A(n2225), .B(n2203), .Z(n1334) );
  CENX1 U2564 ( .A(n2225), .B(n2201), .Z(n1336) );
  CNR2IXL U2565 ( .B(net33082), .A(n2185), .Z(n1054) );
  CENX1 U2566 ( .A(n2238), .B(n2208), .Z(n1268) );
  CENX1 U2567 ( .A(n2228), .B(n2210), .Z(n1326) );
  CENX1 U2568 ( .A(n2240), .B(net33480), .Z(n1277) );
  CENX1 U2569 ( .A(n2242), .B(n1396), .Z(n1270) );
  CENX1 U2570 ( .A(n2246), .B(n2204), .Z(n1246) );
  CENX1 U2571 ( .A(n2246), .B(n2203), .Z(n1247) );
  CENX1 U2572 ( .A(n2246), .B(n2202), .Z(n1248) );
  CENX1 U2573 ( .A(n2239), .B(n2204), .Z(n1273) );
  CENX1 U2574 ( .A(n2240), .B(n2203), .Z(n1274) );
  CENX1 U2575 ( .A(n2246), .B(n2205), .Z(n1245) );
  CENX1 U2576 ( .A(n2238), .B(n2207), .Z(n1269) );
  CENX1 U2577 ( .A(n2238), .B(n2209), .Z(n1267) );
  CENX1 U2578 ( .A(n2248), .B(n2207), .Z(n1242) );
  CENX1 U2579 ( .A(n2241), .B(n2211), .Z(n1265) );
  CENX1 U2580 ( .A(n2235), .B(n2211), .Z(n1294) );
  CENX1 U2581 ( .A(n2241), .B(n2210), .Z(n1266) );
  CENX1 U2582 ( .A(n2248), .B(n2209), .Z(n1240) );
  CENX1 U2583 ( .A(n2206), .B(n2255), .Z(n1196) );
  CENX1 U2584 ( .A(n1396), .B(n2255), .Z(n1195) );
  CENX1 U2585 ( .A(n2241), .B(n2212), .Z(n1264) );
  CENX1 U2586 ( .A(n2208), .B(n2255), .Z(n1193) );
  CENX1 U2587 ( .A(n2207), .B(n2255), .Z(n1194) );
  CENX1 U2588 ( .A(n2209), .B(n2255), .Z(n1192) );
  CENX1 U2589 ( .A(net33482), .B(n2255), .Z(n1203) );
  CENX1 U2590 ( .A(n2219), .B(n2205), .Z(n1365) );
  CENX1 U2591 ( .A(n2205), .B(n2255), .Z(n1197) );
  CENX1 U2592 ( .A(n2225), .B(net33480), .Z(n1337) );
  CENX1 U2593 ( .A(n2228), .B(n2211), .Z(n1325) );
  CENX1 U2594 ( .A(n2226), .B(n2208), .Z(n1328) );
  CENX1 U2595 ( .A(n2228), .B(n2209), .Z(n1327) );
  CENX1 U2596 ( .A(n2235), .B(n2210), .Z(n1295) );
  CENX1 U2597 ( .A(n2226), .B(net33482), .Z(n1338) );
  CENX1 U2598 ( .A(n2235), .B(n2208), .Z(n1297) );
  CENX1 U2599 ( .A(n2234), .B(n2206), .Z(n1300) );
  CENX1 U2600 ( .A(net33082), .B(n2255), .Z(n1204) );
  CENX1 U2601 ( .A(n2224), .B(n2205), .Z(n1332) );
  CENX1 U2602 ( .A(n2224), .B(n2204), .Z(n1333) );
  CENX1 U2603 ( .A(n2228), .B(n2212), .Z(n1324) );
  CNR2X1 U2604 ( .A(n638), .B(n655), .Z(n238) );
  CENX1 U2605 ( .A(net33082), .B(n2235), .Z(n1308) );
  CIVX2 U2606 ( .A(n2237), .Z(n2233) );
  CIVX2 U2607 ( .A(n2237), .Z(n2235) );
  COR2X1 U2608 ( .A(n2025), .B(n2026), .Z(n1035) );
  CNR2XL U2609 ( .A(n18), .B(n1321), .Z(n2025) );
  CNR2XL U2610 ( .A(n1320), .B(n2185), .Z(n2026) );
  CNR2X1 U2611 ( .A(n620), .B(n637), .Z(n233) );
  CND2X1 U2612 ( .A(n638), .B(n655), .Z(n239) );
  CNR2IXL U2613 ( .B(net33082), .A(n1805), .Z(n826) );
  CNR2IXL U2614 ( .B(net33082), .A(n110), .Z(n820) );
  CND2X1 U2615 ( .A(n620), .B(n637), .Z(n234) );
  CND2X1 U2616 ( .A(n2028), .B(n348), .Z(n247) );
  COND2XL U2617 ( .A(n44), .B(n1234), .C(n1233), .D(n42), .Z(n951) );
  CENX1 U2618 ( .A(n246), .B(n132), .Z(product[18]) );
  COND1XL U2619 ( .A(n247), .B(n260), .C(n248), .Z(n246) );
  CND2X1 U2620 ( .A(n346), .B(n245), .Z(n132) );
  CNR2IXL U2621 ( .B(net33082), .A(n6), .Z(product[0]) );
  CENX1 U2622 ( .A(n2248), .B(n1386), .Z(n1233) );
  CENX1 U2623 ( .A(n2229), .B(n1388), .Z(n1322) );
  CENX1 U2624 ( .A(n2223), .B(n1383), .Z(n1317) );
  CENX1 U2625 ( .A(n2223), .B(n1382), .Z(n1316) );
  CENX1 U2626 ( .A(n2238), .B(n1386), .Z(n1260) );
  CENX1 U2627 ( .A(n2231), .B(n1384), .Z(n1287) );
  CENX1 U2628 ( .A(n2223), .B(b[24]), .Z(n1315) );
  CENX1 U2629 ( .A(n2223), .B(b[25]), .Z(n1314) );
  CENX1 U2630 ( .A(n2248), .B(n1385), .Z(n1232) );
  CENX1 U2631 ( .A(n2248), .B(n1384), .Z(n1231) );
  CENX1 U2632 ( .A(n2238), .B(b[24]), .Z(n1255) );
  CENX1 U2633 ( .A(n2238), .B(n1382), .Z(n1256) );
  CENX1 U2634 ( .A(n2238), .B(n1383), .Z(n1257) );
  CENX1 U2635 ( .A(n2248), .B(n1389), .Z(n1236) );
  CENX1 U2636 ( .A(n2248), .B(n1388), .Z(n1235) );
  CENX1 U2637 ( .A(n2248), .B(n1383), .Z(n1230) );
  CENX1 U2638 ( .A(n2236), .B(n1389), .Z(n1292) );
  CENX1 U2639 ( .A(n2236), .B(n1387), .Z(n1290) );
  CENX1 U2640 ( .A(n2231), .B(b[24]), .Z(n1284) );
  CENX1 U2641 ( .A(n2223), .B(b[26]), .Z(n1313) );
  CENX1 U2642 ( .A(n2231), .B(n1383), .Z(n1286) );
  CENX1 U2643 ( .A(n2223), .B(n1386), .Z(n1320) );
  CENX1 U2644 ( .A(n2229), .B(n1389), .Z(n1323) );
  CENX1 U2645 ( .A(n2236), .B(n1388), .Z(n1291) );
  CENX1 U2646 ( .A(n2231), .B(n1385), .Z(n1288) );
  CENX1 U2647 ( .A(n2231), .B(n1382), .Z(n1285) );
  CENX1 U2648 ( .A(n2027), .B(n2127), .Z(n546) );
  CNR2X1 U2649 ( .A(n656), .B(n2092), .Z(n244) );
  CENX1 U2650 ( .A(n2231), .B(n1386), .Z(n1289) );
  CENX1 U2651 ( .A(n2223), .B(b[27]), .Z(n1312) );
  CENX1 U2652 ( .A(n2223), .B(b[28]), .Z(n1311) );
  CENX1 U2653 ( .A(n2231), .B(b[25]), .Z(n1283) );
  CENX1 U2654 ( .A(n2231), .B(b[26]), .Z(n1282) );
  CENX1 U2655 ( .A(n2248), .B(n1387), .Z(n1234) );
  CANR1XL U2656 ( .A(n257), .B(n2028), .C(n250), .Z(n248) );
  COND1XL U2657 ( .A(n2161), .B(n262), .C(n263), .Z(n261) );
  CND2X1 U2658 ( .A(n269), .B(n2182), .Z(n262) );
  CANR1XL U2659 ( .A(n2182), .B(n270), .C(n265), .Z(n263) );
  CENX1 U2660 ( .A(n2241), .B(n1389), .Z(n1263) );
  CENX1 U2661 ( .A(n2239), .B(n1385), .Z(n1259) );
  CENX1 U2662 ( .A(n2239), .B(n1384), .Z(n1258) );
  CENX1 U2663 ( .A(n2219), .B(n1386), .Z(n1353) );
  CENX1 U2664 ( .A(n2219), .B(n1385), .Z(n1352) );
  CENX1 U2665 ( .A(n2219), .B(n1384), .Z(n1351) );
  CENX1 U2666 ( .A(n2219), .B(n1383), .Z(n1350) );
  CENX1 U2667 ( .A(n2219), .B(n1382), .Z(n1349) );
  CENX1 U2668 ( .A(n2219), .B(b[26]), .Z(n1346) );
  CENX1 U2669 ( .A(n2219), .B(b[27]), .Z(n1345) );
  CENX1 U2670 ( .A(n2219), .B(b[24]), .Z(n1348) );
  CENX1 U2671 ( .A(n2219), .B(b[25]), .Z(n1347) );
  CENX1 U2672 ( .A(n2219), .B(b[28]), .Z(n1344) );
  CENX1 U2673 ( .A(n2219), .B(b[29]), .Z(n1343) );
  CENX1 U2674 ( .A(n2219), .B(b[30]), .Z(n1342) );
  CENX1 U2675 ( .A(n2224), .B(n1385), .Z(n1319) );
  CENX1 U2676 ( .A(n2224), .B(n1384), .Z(n1318) );
  COND1XL U2677 ( .A(n2175), .B(n2178), .C(n2177), .Z(n270) );
  CENX1 U2678 ( .A(n2233), .B(b[27]), .Z(n1281) );
  CNR2X1 U2679 ( .A(n2178), .B(n2176), .Z(n269) );
  COR2X1 U2680 ( .A(n2091), .B(n2089), .Z(n2028) );
  CND2X1 U2681 ( .A(n656), .B(n2092), .Z(n245) );
  CEO3X1 U2682 ( .A(n393), .B(n2030), .C(n2031), .Z(n368) );
  CEN3X2 U2683 ( .A(n2155), .B(n403), .C(n2157), .Z(n2030) );
  CEN3X2 U2684 ( .A(n2172), .B(n401), .C(n2159), .Z(n2031) );
  CNIVX2 U2685 ( .A(n1395), .Z(n2207) );
  CNIVX2 U2686 ( .A(n1394), .Z(n2208) );
  CENX1 U2687 ( .A(n2252), .B(n1384), .Z(n1206) );
  CENX1 U2688 ( .A(n2252), .B(n1386), .Z(n1208) );
  CENX1 U2689 ( .A(n2252), .B(n1387), .Z(n1209) );
  CENX1 U2690 ( .A(n2247), .B(n1382), .Z(n1229) );
  CENX1 U2691 ( .A(n2168), .B(n2174), .Z(n2258) );
  CENX1 U2692 ( .A(n278), .B(n137), .Z(product[13]) );
  CND2X1 U2693 ( .A(n351), .B(n2175), .Z(n137) );
  CENX1 U2694 ( .A(n253), .B(n133), .Z(product[17]) );
  COND1XL U2695 ( .A(n2181), .B(n260), .C(n1632), .Z(n253) );
  CENX1 U2696 ( .A(n2226), .B(b[29]), .Z(n1310) );
  CEOX1 U2697 ( .A(n2167), .B(n2173), .Z(n2259) );
  CEOX1 U2698 ( .A(n136), .B(n273), .Z(product[14]) );
  CANR1XL U2699 ( .A(n351), .B(n278), .C(n275), .Z(n273) );
  CEOX1 U2700 ( .A(n135), .B(n268), .Z(n2257) );
  CEOX1 U2701 ( .A(n134), .B(n260), .Z(product[16]) );
  CIVXL U2702 ( .A(n206), .Z(n208) );
  COND2XL U2703 ( .A(n27), .B(n1282), .C(n1281), .D(n2009), .Z(n997) );
  COND2XL U2704 ( .A(n27), .B(n1283), .C(n1282), .D(n2009), .Z(n998) );
  COND2XL U2705 ( .A(n27), .B(n1304), .C(n1303), .D(n2009), .Z(n1019) );
  COND2XL U2706 ( .A(n27), .B(n1301), .C(n1300), .D(n2009), .Z(n1016) );
  COND2XL U2707 ( .A(n27), .B(n1306), .C(n1305), .D(n2009), .Z(n1021) );
  COND2XL U2708 ( .A(n27), .B(n1284), .C(n1283), .D(n2009), .Z(n999) );
  COND2XL U2709 ( .A(n1308), .B(n27), .C(n1307), .D(n2009), .Z(n1023) );
  COND2XL U2710 ( .A(n27), .B(n1302), .C(n1301), .D(n2009), .Z(n1017) );
  COND2XL U2711 ( .A(n27), .B(n2237), .C(n2009), .D(n1309), .Z(n812) );
  COND2XL U2712 ( .A(n27), .B(n1298), .C(n1297), .D(n2009), .Z(n1013) );
  COND2XL U2713 ( .A(n27), .B(n1296), .C(n1295), .D(n2009), .Z(n1011) );
  COND2XL U2714 ( .A(n27), .B(n1289), .C(n1288), .D(n2009), .Z(n1004) );
  COND2XL U2715 ( .A(n27), .B(n1292), .C(n1291), .D(n2009), .Z(n1007) );
  COND2XL U2716 ( .A(n27), .B(n1286), .C(n1285), .D(n2009), .Z(n1001) );
  COND2XL U2717 ( .A(n27), .B(n1290), .C(n1289), .D(n2009), .Z(n1005) );
  COND2XL U2718 ( .A(n1623), .B(n1167), .C(n1166), .D(n1607), .Z(n887) );
  COND2XL U2719 ( .A(n1623), .B(n1169), .C(n1168), .D(n1607), .Z(n889) );
  COND2XL U2720 ( .A(n1623), .B(n1168), .C(n1167), .D(n1607), .Z(n888) );
  COND2XL U2721 ( .A(n1623), .B(n1170), .C(n1169), .D(n1607), .Z(n890) );
  COND2XL U2722 ( .A(n1623), .B(n1171), .C(n1607), .D(n1170), .Z(n891) );
  COND2XL U2723 ( .A(n1623), .B(n1176), .C(n1607), .D(n1175), .Z(n896) );
  COND2XL U2724 ( .A(n1623), .B(n1175), .C(n1607), .D(n1174), .Z(n895) );
  COND2XL U2725 ( .A(n1623), .B(n1177), .C(n1607), .D(n1176), .Z(n897) );
  CND2IXL U2726 ( .B(net33082), .A(n2221), .Z(n1373) );
  COND2XL U2727 ( .A(n1964), .B(n1126), .C(n1555), .D(n1125), .Z(n849) );
  COND2XL U2728 ( .A(n1964), .B(n1131), .C(n89), .D(n1130), .Z(n854) );
  COND2XL U2729 ( .A(n1676), .B(n1122), .C(n1617), .D(n1121), .Z(n845) );
  CND2XL U2730 ( .A(n1035), .B(n981), .Z(n2187) );
  CND2XL U2731 ( .A(n1035), .B(n855), .Z(n2188) );
  CND2XL U2732 ( .A(n981), .B(n855), .Z(n2189) );
  CFA1XL U2733 ( .A(n937), .B(n1067), .CI(n1009), .CO(n649), .S(n650) );
  CND2X1 U2734 ( .A(n565), .B(n546), .Z(n2197) );
  CND2IXL U2735 ( .B(net33082), .A(n1975), .Z(n1228) );
  CIVX2 U2736 ( .A(n2250), .Z(n2246) );
  CND2IXL U2737 ( .B(net33082), .A(n1969), .Z(n1165) );
  CND2IXL U2738 ( .B(net33082), .A(n2215), .Z(n1148) );
  CIVX2 U2739 ( .A(n2230), .Z(n2229) );
  CIVXL U2740 ( .A(n233), .Z(n344) );
  CNR2X1 U2741 ( .A(n233), .B(n238), .Z(n231) );
  CIVX1 U2742 ( .A(n205), .Z(n207) );
  CANR1XL U2743 ( .A(n269), .B(n278), .C(n270), .Z(n268) );
  CND2IXL U2744 ( .B(net33082), .A(n2213), .Z(n1184) );
  CND2X1 U2745 ( .A(n536), .B(n557), .Z(n203) );
  CND2XL U2746 ( .A(n2015), .B(n203), .Z(n126) );
  CND2XL U2747 ( .A(n1844), .B(n214), .Z(n127) );
  CND2X1 U2748 ( .A(n544), .B(n565), .Z(n2195) );
  COND2X1 U2749 ( .A(n53), .B(n1217), .C(n1216), .D(n50), .Z(n935) );
  COND2XL U2750 ( .A(n18), .B(n1311), .C(n1310), .D(n2185), .Z(n1025) );
  COND2XL U2751 ( .A(n18), .B(n1312), .C(n1311), .D(n2185), .Z(n1026) );
  COND2XL U2752 ( .A(n1339), .B(n18), .C(n1338), .D(n2185), .Z(n1053) );
  COND2XL U2753 ( .A(n18), .B(n1337), .C(n1336), .D(n2185), .Z(n1051) );
  COND2XL U2754 ( .A(n18), .B(n1313), .C(n1312), .D(n2185), .Z(n1027) );
  COND2XL U2755 ( .A(n18), .B(n1334), .C(n1333), .D(n2185), .Z(n1048) );
  COND2XL U2756 ( .A(n18), .B(n1325), .C(n1324), .D(n2185), .Z(n1039) );
  COND2XL U2757 ( .A(n18), .B(n1319), .C(n1318), .D(n2185), .Z(n1033) );
  COND2XL U2758 ( .A(n18), .B(n1324), .C(n1323), .D(n2185), .Z(n1038) );
  COND2XL U2759 ( .A(n18), .B(n1328), .C(n1327), .D(n2185), .Z(n1042) );
  CND2XL U2760 ( .A(n538), .B(n559), .Z(n2198) );
  CND2XL U2761 ( .A(n538), .B(n540), .Z(n2199) );
  CND2XL U2762 ( .A(n559), .B(n540), .Z(n2200) );
  CND2X1 U2763 ( .A(n512), .B(n535), .Z(n194) );
  CENX1 U2764 ( .A(n2235), .B(n2209), .Z(n1296) );
  CND2IXL U2765 ( .B(net33082), .A(n2235), .Z(n1309) );
  COND2XL U2766 ( .A(n18), .B(n2230), .C(n2185), .D(n1340), .Z(n813) );
  CND2IXL U2767 ( .B(net33082), .A(n2225), .Z(n1340) );
  COND2XL U2768 ( .A(n44), .B(n2251), .C(n42), .D(n1253), .Z(n810) );
  CND2IXL U2769 ( .B(net33082), .A(n2246), .Z(n1253) );
  CENX1 U2770 ( .A(n2246), .B(n2206), .Z(n1244) );
  CENX1 U2771 ( .A(n2248), .B(n2208), .Z(n1241) );
  CENX1 U2772 ( .A(n2248), .B(n2211), .Z(n1238) );
  CENX1 U2773 ( .A(n2246), .B(n1396), .Z(n1243) );
  CIVX2 U2774 ( .A(n2245), .Z(n2241) );
  COND2XL U2775 ( .A(n9), .B(n2222), .C(n6), .D(n1373), .Z(n814) );
  CND2IXL U2776 ( .B(net33082), .A(n2238), .Z(n1280) );
  CEOXL U2777 ( .A(n309), .B(n143), .Z(product[7]) );
  CEOXL U2778 ( .A(n317), .B(n145), .Z(product[5]) );
  COND1XL U2779 ( .A(n205), .B(n222), .C(n1903), .Z(n204) );
  COND2XL U2780 ( .A(n53), .B(n1207), .C(n1206), .D(n50), .Z(n925) );
  COND2XL U2781 ( .A(n53), .B(n1208), .C(n1207), .D(n50), .Z(n926) );
  COND2XL U2782 ( .A(n53), .B(n1209), .C(n1208), .D(n50), .Z(n927) );
  COND2XL U2783 ( .A(n53), .B(n1211), .C(n1210), .D(n50), .Z(n929) );
  COND2XL U2784 ( .A(n53), .B(n1210), .C(n1209), .D(n50), .Z(n928) );
  COND2XL U2785 ( .A(n53), .B(n1220), .C(n1219), .D(n50), .Z(n938) );
  COND2XL U2786 ( .A(n53), .B(n1221), .C(n1220), .D(n50), .Z(n939) );
  COND2XL U2787 ( .A(n53), .B(n1219), .C(n1218), .D(n50), .Z(n937) );
  COND2XL U2788 ( .A(n53), .B(n1225), .C(n1224), .D(n50), .Z(n943) );
  COND2XL U2789 ( .A(n53), .B(n1213), .C(n1212), .D(n50), .Z(n931) );
  COND2XL U2790 ( .A(n53), .B(n1216), .C(n1215), .D(n50), .Z(n934) );
  COND2XL U2791 ( .A(n53), .B(n1215), .C(n1214), .D(n50), .Z(n933) );
  COND2XL U2792 ( .A(n53), .B(n1212), .C(n1211), .D(n50), .Z(n930) );
  COND2XL U2793 ( .A(n53), .B(n1222), .C(n1221), .D(n50), .Z(n940) );
  COND2XL U2794 ( .A(n53), .B(n1214), .C(n1213), .D(n50), .Z(n932) );
  COND2XL U2795 ( .A(n53), .B(n1218), .C(n1217), .D(n50), .Z(n936) );
  CIVX4 U2796 ( .A(a[0]), .Z(n6) );
  CND2X4 U2797 ( .A(n1421), .B(n6), .Z(n9) );
  CND2X4 U2798 ( .A(n1420), .B(n2184), .Z(n18) );
  CND2X4 U2799 ( .A(n1418), .B(n33), .Z(n36) );
  CND2X4 U2800 ( .A(n1417), .B(n42), .Z(n44) );
  CIVXL U2801 ( .A(n2230), .Z(n2223) );
  CIVXL U2802 ( .A(n2237), .Z(n2231) );
  CIVXL U2803 ( .A(n2237), .Z(n2232) );
  CIVXL U2804 ( .A(n2237), .Z(n2236) );
  CIVXL U2805 ( .A(n30), .Z(n2243) );
  CIVXL U2806 ( .A(n2251), .Z(n2249) );
  CIVX2 U2807 ( .A(n323), .Z(n361) );
  CIVX2 U2808 ( .A(n2178), .Z(n350) );
  CIVX2 U2809 ( .A(n244), .Z(n346) );
  CIVX2 U2810 ( .A(n332), .Z(n330) );
  CIVX2 U2811 ( .A(n329), .Z(n327) );
  CIVX2 U2812 ( .A(n321), .Z(n319) );
  CIVX2 U2813 ( .A(n313), .Z(n311) );
  CIVX2 U2814 ( .A(n305), .Z(n303) );
  CIVX2 U2815 ( .A(n2175), .Z(n275) );
  CIVX2 U2816 ( .A(n2176), .Z(n351) );
  CIVX2 U2817 ( .A(n2179), .Z(n265) );
  CIVX2 U2818 ( .A(n2180), .Z(n257) );
  CIVX2 U2819 ( .A(n2181), .Z(n348) );
  CIVX2 U2820 ( .A(n252), .Z(n250) );
  CIVX2 U2821 ( .A(n241), .Z(n240) );
  CIVX2 U2822 ( .A(n239), .Z(n237) );
  CIVX2 U2823 ( .A(n238), .Z(n345) );
  CIVX2 U2824 ( .A(n217), .Z(n219) );
  CIVX2 U2825 ( .A(n216), .Z(n342) );
  CIVX2 U2826 ( .A(n203), .Z(n201) );
endmodule


module calc_DW02_mult_2_stage_0 ( A, B, TC, CLK, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC, CLK;
  wire   n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         \A_extended[32] , \B_extended[32] , n6, n8, n10, n12, n14, n16, n18,
         n19, n21, n23, n25, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33;
  assign \A_extended[32]  = A[31];
  assign \B_extended[32]  = B[31];

  calc_DW_mult_tc_23 mult_96 ( .a({\A_extended[32] , \A_extended[32] , A[30:0]}), .b({\B_extended[32] , \B_extended[32] , B[30:0]}), .product({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, PRODUCT[31:12], 
        n39, PRODUCT[10], n40, n41, n42, n43, n44, n45, n46, n47, n48, n49}), 
        .i_retiming_group_0_clk(CLK) );
  CFD1QXL clk_r_REG166_S1 ( .D(n49), .CP(CLK), .Q(n28) );
  CFD1QXL clk_r_REG136_S1 ( .D(n48), .CP(CLK), .Q(n29) );
  CFD1QXL clk_r_REG77_S1 ( .D(n43), .CP(CLK), .Q(n34) );
  CFD1QXL clk_r_REG86_S1 ( .D(n44), .CP(CLK), .Q(n33) );
  CFD1QXL clk_r_REG90_S1 ( .D(n45), .CP(CLK), .Q(n32) );
  CFD1QXL clk_r_REG100_S1 ( .D(n46), .CP(CLK), .Q(n31) );
  CFD1QXL clk_r_REG104_S1 ( .D(n47), .CP(CLK), .Q(n30) );
  CFD1QXL clk_r_REG0_S1 ( .D(n40), .CP(CLK), .Q(n37) );
  CFD1QXL clk_r_REG56_S1 ( .D(n41), .CP(CLK), .Q(n36) );
  CFD1QX2 clk_r_REG3_S1 ( .D(n39), .CP(CLK), .Q(n38) );
  CFD1QXL clk_r_REG63_S1 ( .D(n42), .CP(CLK), .Q(n35) );
  CIVDXL U1 ( .A(n37), .Z1(n6) );
  CNIVX1 U2 ( .A(n6), .Z(PRODUCT[9]) );
  CIVDXL U3 ( .A(n34), .Z1(n8) );
  CNIVX1 U4 ( .A(n8), .Z(PRODUCT[6]) );
  CIVDXL U5 ( .A(n30), .Z1(n10) );
  CNIVX1 U6 ( .A(n10), .Z(PRODUCT[2]) );
  CIVDXL U7 ( .A(n36), .Z1(n12) );
  CNIVX1 U8 ( .A(n12), .Z(PRODUCT[8]) );
  CIVDXL U9 ( .A(n33), .Z1(n14) );
  CNIVX1 U10 ( .A(n14), .Z(PRODUCT[5]) );
  CIVDXL U11 ( .A(n32), .Z1(n16) );
  CNIVX1 U12 ( .A(n16), .Z(PRODUCT[4]) );
  CNIVX3 U13 ( .A(n38), .Z(n19) );
  CNIVX1 U14 ( .A(n18), .Z(PRODUCT[11]) );
  CNIVX1 U15 ( .A(n19), .Z(n18) );
  CIVDXL U16 ( .A(n31), .Z1(n21) );
  CNIVX1 U17 ( .A(n21), .Z(PRODUCT[3]) );
  CIVDXL U18 ( .A(n28), .Z1(n23) );
  CNIVX1 U19 ( .A(n23), .Z(PRODUCT[0]) );
  CIVDXL U20 ( .A(n35), .Z1(n25) );
  CNIVX1 U21 ( .A(n25), .Z(PRODUCT[7]) );
  CIVDXL U22 ( .A(n29), .Z1(n27) );
  CNIVX1 U23 ( .A(n27), .Z(PRODUCT[1]) );
endmodule


module calc_DW_mult_tc_22 ( a, b, product, i_retiming_group_0_clk );
  input [32:0] a;
  input [32:0] b;
  output [65:0] product;
  input i_retiming_group_0_clk;
  wire   n3, n6, n9, n12, n15, n18, n21, n24, n27, n30, n36, n39, n42, n44,
         n48, n50, n53, n55, n58, n61, n63, n66, n69, n71, n74, n77, n79, n82,
         n84, n86, n89, n91, n93, n95, n97, n99, n100, n102, n104, n105, n107,
         n109, n116, n119, n120, n123, n124, n125, n127, n129, n131, n132,
         n133, n136, n137, n138, n139, n141, n142, n143, n144, n145, n146,
         n147, n148, n151, n154, n156, n157, n158, n159, n160, n161, n163,
         n164, n165, n166, n167, n170, n171, n172, n173, n175, n178, n179,
         n182, n183, n184, n185, n195, n196, n197, n205, n208, n215, n216,
         n222, n229, n230, n231, n232, n233, n234, n235, n237, n238, n239,
         n244, n245, n246, n247, n248, n251, n252, n253, n254, n255, n260,
         n261, n262, n263, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n288, n289, n290, n292, n294, n295, n297, n299, n300,
         n301, n303, n305, n306, n307, n308, n309, n311, n313, n314, n315,
         n316, n317, n319, n321, n322, n323, n324, n325, n327, n329, n330,
         n332, n335, n336, n337, n342, n344, n345, n346, n347, n348, n349,
         n351, n353, n361, n364, n365, n368, n369, n370, n371, n372, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n427, n429, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n541, n542, n543, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n558, n560, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n820, n821, n822, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1089, n1090, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1408, n1409, n1411, n1412, n1415,
         n1416, n1418, n1420, n1421, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, net32098, net33078, net33076, net33422, net33757,
         net33755, net33754, net33752, net171472, net171496, net171498,
         net171589, net171591, net171592, net171593, net171594, net171595,
         net171596, net171597, net171598, net171599, net171600, net171602,
         net171604, net171605, net178512, net178605, net178660, net178746,
         net178962, net179383, net179382, net179418, net179429, net179428,
         net179427, net179529, net179547, net179546, net179617, net179825,
         net179824, net179820, net179838, net179858, net179943, net179942,
         net179941, net180011, net180068, net180217, net180366, net180365,
         net180364, net180562, net180674, net180673, net181698, net179676,
         n243, n242, n227, n225, n224, n223, n186, net33776, net33775,
         net33774, net180618, net180312, net179842, net178513, net178507, n579,
         n512, n217, n214, n212, n206, n194, n192, n190, n189, n188, n187,
         n566, net182741, n799, n1088, n1087, n1086, net183987, net184278,
         net184277, net184424, n1091, net183988, net182674, net182673,
         net182672, n1407, n112, n110, net184434, net184082, n973, n907, n823,
         n819, n430, n428, n426, n1092, n1057, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205;
  assign n3 = a[1];
  assign n12 = a[3];
  assign n21 = a[5];
  assign n30 = a[7];
  assign n39 = a[9];
  assign n48 = a[11];
  assign n55 = a[13];
  assign n63 = a[15];
  assign n71 = a[17];
  assign n79 = a[19];
  assign n86 = a[21];
  assign n93 = a[23];
  assign n99 = a[25];
  assign n104 = a[27];
  assign n109 = a[29];
  assign n116 = b[0];
  assign n1382 = b[23];
  assign n1383 = b[22];
  assign n1384 = b[21];
  assign n1385 = b[20];
  assign n1386 = b[19];
  assign n1387 = b[18];
  assign n1388 = b[17];
  assign n1389 = b[16];
  assign n1390 = b[15];
  assign n1391 = b[14];
  assign n1392 = b[13];
  assign n1393 = b[12];
  assign n1394 = b[11];
  assign n1395 = b[10];
  assign n1396 = b[9];
  assign n1397 = b[8];
  assign n1398 = b[7];
  assign n1399 = b[6];
  assign n1400 = b[5];
  assign n1401 = b[4];
  assign n1402 = b[3];
  assign n1403 = b[2];
  assign n1404 = b[1];
  assign n2114 = i_retiming_group_0_clk;

  CANR1X1 U119 ( .A(n165), .B(n185), .C(n1636), .Z(n164) );
  CNR2X2 U214 ( .A(n620), .B(n637), .Z(n233) );
  CANR1X1 U217 ( .A(n345), .B(n1662), .C(n237), .Z(n235) );
  CEO3X2 U371 ( .A(n383), .B(n365), .C(n381), .Z(n364) );
  CEO3X2 U375 ( .A(n2091), .B(n2098), .C(n2099), .Z(n368) );
  CFA1X1 U386 ( .A(n384), .B(n382), .CI(n409), .CO(n379), .S(n380) );
  CFA1X1 U387 ( .A(n388), .B(n411), .CI(n386), .CO(n381), .S(n382) );
  CFA1X1 U388 ( .A(n2094), .B(n413), .CI(n415), .CO(n383), .S(n384) );
  CFA1X1 U389 ( .A(n2088), .B(n2092), .CI(n2090), .CO(n385), .S(n386) );
  CFA1X1 U390 ( .A(n2084), .B(n2089), .CI(n2086), .CO(n387), .S(n388) );
  CFA1X1 U395 ( .A(n972), .B(n1056), .CI(n1026), .CO(n397), .S(n398) );
  CFA1X1 U399 ( .A(n1811), .B(n836), .CI(n816), .CO(n405), .S(n406) );
  CFA1X1 U400 ( .A(n412), .B(n410), .CI(n437), .CO(n407), .S(n408) );
  CFA1X1 U401 ( .A(n416), .B(n439), .CI(n414), .CO(n409), .S(n410) );
  CFA1X1 U402 ( .A(n2087), .B(n441), .CI(n443), .CO(n411), .S(n412) );
  CFA1X1 U403 ( .A(n2083), .B(n2085), .CI(n2081), .CO(n413), .S(n414) );
  CFA1X1 U404 ( .A(n2077), .B(n2079), .CI(n2082), .CO(n415), .S(n416) );
  CFA1X1 U407 ( .A(n457), .B(n455), .CI(n459), .CO(n421), .S(n422) );
  CFA1X1 U408 ( .A(n999), .B(n434), .CI(n1027), .CO(n423), .S(n424) );
  CFA1X1 U417 ( .A(n2076), .B(n2078), .CI(n2074), .CO(n441), .S(n442) );
  CFA1X1 U418 ( .A(n2075), .B(n2072), .CI(n2070), .CO(n443), .S(n444) );
  CFA1X1 U422 ( .A(n1000), .B(n1058), .CI(n1028), .CO(n451), .S(n452) );
  CFA1X1 U427 ( .A(n466), .B(n464), .CI(n489), .CO(n461), .S(n462) );
  CFA1X1 U428 ( .A(n470), .B(n491), .CI(n468), .CO(n463), .S(n464) );
  CFA1X1 U432 ( .A(n484), .B(n480), .CI(n501), .CO(n471), .S(n472) );
  CFA1X1 U433 ( .A(n505), .B(n503), .CI(n507), .CO(n473), .S(n474) );
  CFA1X1 U434 ( .A(n1029), .B(n509), .CI(n486), .CO(n475), .S(n476) );
  CFA1X1 U435 ( .A(n1001), .B(n825), .CI(n1059), .CO(n477), .S(n478) );
  CHA1X1 U439 ( .A(n849), .B(n891), .CO(n485), .S(n486) );
  CFA1X1 U440 ( .A(n492), .B(n513), .CI(n490), .CO(n487), .S(n488) );
  CFA1X1 U441 ( .A(n517), .B(n515), .CI(n494), .CO(n489), .S(n490) );
  CFA1X1 U442 ( .A(n2060), .B(n2065), .CI(n2063), .CO(n491), .S(n492) );
  CFA1X1 U443 ( .A(n2058), .B(n2061), .CI(n2096), .CO(n493), .S(n494) );
  CFA1X1 U444 ( .A(n502), .B(n506), .CI(n504), .CO(n495), .S(n496) );
  CFA1X1 U445 ( .A(n525), .B(n508), .CI(n510), .CO(n497), .S(n498) );
  CFA1X1 U446 ( .A(n531), .B(n527), .CI(n529), .CO(n499), .S(n500) );
  CFA1X1 U447 ( .A(n1002), .B(n533), .CI(n1030), .CO(n501), .S(n502) );
  CFA1X1 U454 ( .A(n2059), .B(n543), .CI(n2102), .CO(n515), .S(n516) );
  CFA1X1 U455 ( .A(n2055), .B(n2057), .CI(n2056), .CO(n517), .S(n518) );
  CFA1X1 U456 ( .A(n528), .B(n530), .CI(n526), .CO(n519), .S(n520) );
  CFA1X1 U460 ( .A(n911), .B(n1061), .CI(n977), .CO(n527), .S(n528) );
  CHA1X1 U463 ( .A(n863), .B(n893), .CO(n533), .S(n534) );
  CFA1X1 U470 ( .A(n1004), .B(n575), .CI(n577), .CO(n547), .S(n548) );
  CFA1X1 U471 ( .A(n978), .B(n1062), .CI(n1032), .CO(n549), .S(n550) );
  CFA1X1 U481 ( .A(n1005), .B(n578), .CI(n1033), .CO(n569), .S(n570) );
  CFA1X1 U487 ( .A(n2053), .B(n2052), .CI(n2054), .CO(n581), .S(n582) );
  CFA1X1 U489 ( .A(n594), .B(n609), .CI(n592), .CO(n585), .S(n586) );
  CFA1X1 U490 ( .A(n611), .B(n596), .CI(n598), .CO(n587), .S(n588) );
  CFA1X1 U492 ( .A(n980), .B(n1034), .CI(n1006), .CO(n591), .S(n592) );
  CFA1X1 U502 ( .A(n981), .B(n855), .CI(n1035), .CO(n611), .S(n612) );
  CFA1X1 U507 ( .A(n2046), .B(n2043), .CI(n2103), .CO(n621), .S(n622) );
  CFA1X1 U508 ( .A(n630), .B(n643), .CI(n645), .CO(n623), .S(n624) );
  CFA1X1 U510 ( .A(n651), .B(n649), .CI(n647), .CO(n627), .S(n628) );
  CFA1X1 U511 ( .A(n958), .B(n653), .CI(n982), .CO(n629), .S(n630) );
  CFA1X1 U515 ( .A(n2042), .B(n2044), .CI(n2041), .CO(n637), .S(n638) );
  CFA1X1 U516 ( .A(n646), .B(n644), .CI(n659), .CO(n639), .S(n640) );
  CFA1X1 U517 ( .A(n648), .B(n661), .CI(n663), .CO(n641), .S(n642) );
  CFA1X1 U520 ( .A(n959), .B(n869), .CI(n983), .CO(n647), .S(n648) );
  CFA1X1 U522 ( .A(n1967), .B(n805), .CI(n1037), .CO(n651), .S(n652) );
  CHA1X1 U523 ( .A(n917), .B(n883), .CO(n653), .S(n654) );
  CFA1X1 U526 ( .A(n666), .B(n677), .CI(n679), .CO(n659), .S(n660) );
  CFA1X1 U528 ( .A(n984), .B(n683), .CI(n685), .CO(n663), .S(n664) );
  CFA1X1 U531 ( .A(n870), .B(n884), .CI(n1965), .CO(n669), .S(n670) );
  CFA1X1 U532 ( .A(n2037), .B(n2036), .CI(n2033), .CO(n671), .S(n672) );
  CFA1X1 U533 ( .A(n680), .B(n691), .CI(n678), .CO(n673), .S(n674) );
  CFA1X1 U534 ( .A(n684), .B(n693), .CI(n682), .CO(n675), .S(n676) );
  CFA1X1 U535 ( .A(n695), .B(n699), .CI(n697), .CO(n677), .S(n678) );
  CFA1X1 U536 ( .A(n1011), .B(n686), .CI(n1039), .CO(n679), .S(n680) );
  CFA1X1 U537 ( .A(n919), .B(n885), .CI(n985), .CO(n681), .S(n682) );
  CFA1X1 U540 ( .A(n692), .B(n690), .CI(n703), .CO(n687), .S(n688) );
  CFA1X1 U541 ( .A(n707), .B(n694), .CI(n705), .CO(n689), .S(n690) );
  CFA1X1 U542 ( .A(n696), .B(n700), .CI(n698), .CO(n691), .S(n692) );
  CFA1X1 U543 ( .A(n711), .B(n709), .CI(n713), .CO(n693), .S(n694) );
  CFA1X1 U544 ( .A(n962), .B(n1040), .CI(n986), .CO(n695), .S(n696) );
  CFA1X1 U554 ( .A(n720), .B(n718), .CI(n729), .CO(n715), .S(n716) );
  CFA1X1 U555 ( .A(n724), .B(n731), .CI(n722), .CO(n717), .S(n718) );
  CFA1X1 U557 ( .A(n988), .B(n737), .CI(n1014), .CO(n721), .S(n722) );
  CFA1X1 U560 ( .A(n732), .B(n730), .CI(n741), .CO(n727), .S(n728) );
  CFA1X1 U561 ( .A(n736), .B(n734), .CI(n743), .CO(n729), .S(n730) );
  CFA1X1 U562 ( .A(n738), .B(n745), .CI(n747), .CO(n731), .S(n732) );
  CFA1X1 U566 ( .A(n751), .B(n742), .CI(n744), .CO(n739), .S(n740) );
  CFA1X1 U567 ( .A(n748), .B(n753), .CI(n746), .CO(n741), .S(n742) );
  CFA1X1 U568 ( .A(n1016), .B(n755), .CI(n757), .CO(n743), .S(n744) );
  CFA1X1 U571 ( .A(n754), .B(n752), .CI(n761), .CO(n749), .S(n750) );
  CFA1X1 U572 ( .A(n765), .B(n756), .CI(n763), .CO(n751), .S(n752) );
  CFA1X1 U573 ( .A(n991), .B(n758), .CI(n1017), .CO(n753), .S(n754) );
  CFA1X1 U574 ( .A(n967), .B(n1075), .CI(n1045), .CO(n755), .S(n756) );
  CFA1X1 U576 ( .A(n764), .B(n762), .CI(n769), .CO(n759), .S(n760) );
  CFA1X1 U577 ( .A(n773), .B(n766), .CI(n771), .CO(n761), .S(n762) );
  CFA1X1 U578 ( .A(n1018), .B(n1076), .CI(n1046), .CO(n763), .S(n764) );
  CFA1X1 U580 ( .A(n777), .B(n770), .CI(n772), .CO(n767), .S(n768) );
  CFA1X1 U581 ( .A(n1019), .B(n779), .CI(n774), .CO(n769), .S(n770) );
  CFA1X1 U582 ( .A(n1665), .B(n969), .CI(n1047), .CO(n771), .S(n772) );
  CHA1X1 U583 ( .A(n810), .B(n1077), .CO(n773), .S(n774) );
  CFA1X1 U584 ( .A(n783), .B(n778), .CI(n780), .CO(n775), .S(n776) );
  CFA1X1 U585 ( .A(n1048), .B(n785), .CI(n1078), .CO(n777), .S(n778) );
  CFA1X1 U586 ( .A(n970), .B(n1020), .CI(n994), .CO(n779), .S(n780) );
  CFA1X1 U587 ( .A(n786), .B(n784), .CI(n789), .CO(n781), .S(n782) );
  CFA1X1 U588 ( .A(n1021), .B(n1079), .CI(n1667), .CO(n783), .S(n784) );
  CHA1X1 U589 ( .A(n811), .B(n995), .CO(n785), .S(n786) );
  CFA1X1 U592 ( .A(n1051), .B(n794), .CI(n1081), .CO(n791), .S(n792) );
  CHA1X1 U593 ( .A(n812), .B(n1023), .CO(n793), .S(n794) );
  CFA1X1 U594 ( .A(n1024), .B(n1082), .CI(n1052), .CO(n795), .S(n796) );
  CHA1X1 U595 ( .A(n813), .B(n1083), .CO(n797), .S(n798) );
  COND2X1 U616 ( .A(n107), .B(n1098), .C(net181698), .D(n1097), .Z(n824) );
  COND2X1 U617 ( .A(n107), .B(n1099), .C(net181698), .D(n1098), .Z(n825) );
  COND2X1 U628 ( .A(n1103), .B(n1747), .C(n1814), .D(n1102), .Z(n828) );
  COND2X1 U629 ( .A(n1104), .B(n1747), .C(n1814), .D(n1103), .Z(n829) );
  COND2X1 U633 ( .A(n102), .B(n1108), .C(n1814), .D(n1737), .Z(n833) );
  COND2X1 U704 ( .A(n84), .B(n1146), .C(n82), .D(n1145), .Z(n868) );
  COND2X1 U733 ( .A(n1697), .B(n1160), .C(n74), .D(n1159), .Z(n881) );
  COND2X1 U736 ( .A(n77), .B(n1163), .C(n74), .D(n1162), .Z(n884) );
  COND2X1 U904 ( .A(n44), .B(n1251), .C(n1250), .D(n42), .Z(n968) );
  CND2IX1 U931 ( .B(net33078), .A(n2191), .Z(n1253) );
  COND2X1 U990 ( .A(n27), .B(n1285), .C(n1284), .D(n24), .Z(n1000) );
  COND2X1 U991 ( .A(n27), .B(n1286), .C(n1285), .D(n24), .Z(n1001) );
  COND2X1 U992 ( .A(n27), .B(n1287), .C(n1286), .D(n24), .Z(n1002) );
  COND2X1 U995 ( .A(n27), .B(n1290), .C(n1289), .D(n24), .Z(n1005) );
  COND2X1 U996 ( .A(n27), .B(n1291), .C(n1290), .D(n24), .Z(n1006) );
  COND2X1 U998 ( .A(n27), .B(n1293), .C(n1292), .D(n24), .Z(n1008) );
  COND2X1 U999 ( .A(n27), .B(n1294), .C(n1293), .D(n24), .Z(n1009) );
  COND2X1 U1000 ( .A(n27), .B(n1295), .C(n1294), .D(n24), .Z(n1010) );
  COND2X1 U1002 ( .A(n27), .B(n1297), .C(n1296), .D(n24), .Z(n1012) );
  COND2X1 U1004 ( .A(n27), .B(n1299), .C(n1298), .D(n24), .Z(n1014) );
  COND2X1 U1005 ( .A(n27), .B(n1300), .C(n1299), .D(n24), .Z(n1015) );
  COND2X1 U1010 ( .A(n27), .B(n1305), .C(n1304), .D(n24), .Z(n1020) );
  CND2IX1 U1043 ( .B(net33078), .A(n2176), .Z(n1309) );
  COND2X1 U1047 ( .A(n18), .B(n1313), .C(n1312), .D(n15), .Z(n1027) );
  COND2X1 U1048 ( .A(n18), .B(n1314), .C(n1313), .D(n15), .Z(n1028) );
  COND2X1 U1050 ( .A(n18), .B(n1316), .C(n1315), .D(n15), .Z(n1030) );
  COND2X1 U1052 ( .A(n18), .B(n1318), .C(n1317), .D(n15), .Z(n1032) );
  COND2X1 U1054 ( .A(n18), .B(n1320), .C(n1319), .D(n15), .Z(n1034) );
  COND2X1 U1055 ( .A(n18), .B(n1321), .C(n1320), .D(n15), .Z(n1035) );
  COND2X1 U1057 ( .A(n18), .B(n1323), .C(n1322), .D(n15), .Z(n1037) );
  COND2X1 U1058 ( .A(n18), .B(n1324), .C(n1323), .D(n15), .Z(n1038) );
  COND2X1 U1060 ( .A(n18), .B(n1326), .C(n1325), .D(n15), .Z(n1040) );
  COND2X1 U1062 ( .A(n18), .B(n1328), .C(n1327), .D(n15), .Z(n1042) );
  COND2X1 U1063 ( .A(n18), .B(n1329), .C(n1328), .D(n15), .Z(n1043) );
  COND2X1 U1064 ( .A(n18), .B(n1330), .C(n1329), .D(n15), .Z(n1044) );
  COND2X1 U1065 ( .A(n18), .B(n1331), .C(n1330), .D(n15), .Z(n1045) );
  COND2X1 U1067 ( .A(n18), .B(n1333), .C(n1332), .D(n15), .Z(n1047) );
  COND2X1 U1107 ( .A(n1548), .B(n1342), .C(n6), .D(n1341), .Z(n1055) );
  COND2X1 U1111 ( .A(n1548), .B(n1346), .C(n6), .D(n1345), .Z(n1059) );
  COND2X1 U1112 ( .A(n1548), .B(n1347), .C(n6), .D(n1346), .Z(n1060) );
  COND2X1 U1113 ( .A(n1548), .B(n1348), .C(n6), .D(n1347), .Z(n1061) );
  COND2X1 U1114 ( .A(n1548), .B(n1349), .C(n6), .D(n1348), .Z(n1062) );
  COND2X1 U1115 ( .A(n1548), .B(n1350), .C(n6), .D(n1349), .Z(n1063) );
  COND2X1 U1116 ( .A(n1548), .B(n1351), .C(n6), .D(n1350), .Z(n1064) );
  COND2X1 U1117 ( .A(n1548), .B(n1352), .C(n6), .D(n1351), .Z(n1065) );
  COND2X1 U1118 ( .A(n1548), .B(n1353), .C(n6), .D(n1352), .Z(n1066) );
  COND2X1 U1119 ( .A(n9), .B(n1354), .C(n6), .D(n1353), .Z(n1067) );
  COND2X1 U1120 ( .A(n9), .B(n1355), .C(n6), .D(n1354), .Z(n1068) );
  COND2X1 U1121 ( .A(n1548), .B(n1356), .C(n6), .D(n1355), .Z(n1069) );
  COND2X1 U1122 ( .A(n9), .B(n1357), .C(n6), .D(n1356), .Z(n1070) );
  COND2X1 U1123 ( .A(n9), .B(n1358), .C(n6), .D(n1357), .Z(n1071) );
  COND2X1 U1124 ( .A(n9), .B(n1359), .C(n6), .D(n1358), .Z(n1072) );
  COND2X1 U1125 ( .A(n9), .B(n1360), .C(n6), .D(n1359), .Z(n1073) );
  COND2X1 U1126 ( .A(n9), .B(n1361), .C(n6), .D(n1360), .Z(n1074) );
  COND2X1 U1127 ( .A(n9), .B(n1362), .C(n6), .D(n1361), .Z(n1075) );
  COND2X1 U1128 ( .A(n9), .B(n1363), .C(n6), .D(n1362), .Z(n1076) );
  COND2X1 U1129 ( .A(n9), .B(n1364), .C(n6), .D(n1363), .Z(n1077) );
  COND2X1 U1130 ( .A(n9), .B(n1365), .C(n6), .D(n1364), .Z(n1078) );
  COND2X1 U1131 ( .A(n9), .B(n1366), .C(n6), .D(n1365), .Z(n1079) );
  COND2X1 U1132 ( .A(n9), .B(n1367), .C(n6), .D(n1366), .Z(n1080) );
  COND2X1 U1133 ( .A(n9), .B(n1368), .C(n6), .D(n1367), .Z(n1081) );
  COND2X1 U1134 ( .A(n9), .B(n1369), .C(n6), .D(n1368), .Z(n1082) );
  COND2X1 U1135 ( .A(n9), .B(n1370), .C(n6), .D(n1369), .Z(n1083) );
  COND2X1 U1136 ( .A(n9), .B(n1371), .C(n6), .D(n1370), .Z(n1084) );
  COND2X1 U1137 ( .A(n9), .B(n1372), .C(n6), .D(n1371), .Z(n1085) );
  CEOX2 U1254 ( .A(a[6]), .B(n2187), .Z(n1418) );
  CEOX2 U1260 ( .A(a[2]), .B(n2171), .Z(n1420) );
  CFD1QX1 clk_r_REG175_S1 ( .D(n687), .CP(n2114), .Q(n2035) );
  CFD1QX1 clk_r_REG172_S1 ( .D(n701), .CP(n2114), .Q(n2032) );
  CFD1QXL clk_r_REG265_S1 ( .D(n393), .CP(n2114), .Q(n2091) );
  CFD1QXL clk_r_REG272_S1 ( .D(n371), .CP(n2114), .Q(n2099) );
  CFD1QXL clk_r_REG243_S1 ( .D(n396), .CP(n2114), .Q(n2089) );
  CFD1QXL clk_r_REG241_S1 ( .D(n389), .CP(n2114), .Q(n2095) );
  CFD1QXL clk_r_REG239_S1 ( .D(n372), .CP(n2114), .Q(n2098) );
  CFD1QXL clk_r_REG266_S1 ( .D(n394), .CP(n2114), .Q(n2090) );
  CFD1QXL clk_r_REG179_S1 ( .D(n657), .CP(n2114), .Q(n2041) );
  CFD1QXL clk_r_REG184_S1 ( .D(n639), .CP(n2114), .Q(n2045) );
  CFD1QXL clk_r_REG188_S1 ( .D(n421), .CP(n2114), .Q(n2084) );
  CFD1QXL clk_r_REG196_S1 ( .D(n642), .CP(n2114), .Q(n2042) );
  CFD1QXL clk_r_REG198_S1 ( .D(n624), .CP(n2114), .Q(n2047) );
  CFD1QXL clk_r_REG202_S1 ( .D(n138), .CP(n2114), .Q(n2106) );
  CFD1QXL clk_r_REG221_S1 ( .D(n495), .CP(n2114), .Q(n2066) );
  CFD1QX2 clk_r_REG210_S1 ( .D(n554), .CP(n2114), .Q(net171592) );
  CFD1QX2 clk_r_REG235_S1 ( .D(n626), .CP(n2114), .Q(n2103) );
  CFD1QX2 clk_r_REG257_S1 ( .D(n576), .CP(n2114), .Q(net171597) );
  CFD1QX2 clk_r_REG204_S1 ( .D(n276), .CP(n2114), .Q(n2108) );
  CFD1QX2 clk_r_REG280_S1 ( .D(n574), .CP(n2114), .Q(net171596) );
  CFD1QX2 clk_r_REG213_S1 ( .D(n570), .CP(n2114), .Q(net171594) );
  CFD1QX2 clk_r_REG183_S1 ( .D(n660), .CP(n2114), .Q(n2039) );
  CFD1QX1 clk_r_REG195_S1 ( .D(n641), .CP(n2114), .Q(n2043) );
  CFD1QX2 clk_r_REG201_S1 ( .D(n285), .CP(n2114), .Q(n2105) );
  CFD1QX1 clk_r_REG181_S1 ( .D(n673), .CP(n2114), .Q(n2038) );
  CFD1QX2 clk_r_REG245_S1 ( .D(n497), .CP(n2114), .Q(n2064) );
  CFD1QX1 clk_r_REG219_S1 ( .D(n499), .CP(n2114), .Q(n2062) );
  CFD1QX2 clk_r_REG250_S1 ( .D(n587), .CP(n2114), .Q(net171602) );
  CFD1QX2 clk_r_REG187_S1 ( .D(n446), .CP(n2114), .Q(n2080) );
  CFD1QX2 clk_r_REG206_S1 ( .D(n271), .CP(n2114), .Q(n2110) );
  CFD1QX2 clk_r_REG254_S1 ( .D(n448), .CP(n2114), .Q(n2078) );
  CFD1QX2 clk_r_REG224_S1 ( .D(n474), .CP(n2114), .Q(n2071) );
  CFD1QX2 clk_r_REG173_S1 ( .D(n267), .CP(n2114), .Q(n2111) );
  CFD1QX2 clk_r_REG256_S1 ( .D(n420), .CP(n2114), .Q(n2085) );
  CFD1QX1 clk_r_REG197_S1 ( .D(n623), .CP(n2114), .Q(n2048) );
  CFD1QX2 clk_r_REG174_S1 ( .D(n266), .CP(n2114), .Q(n2112) );
  CFD1QX1 clk_r_REG192_S1 ( .D(n449), .CP(n2114), .Q(n2077) );
  CFD1QX2 clk_r_REG231_S1 ( .D(n589), .CP(n2114), .Q(net171604) );
  CFD1QX1 clk_r_REG274_S1 ( .D(n452), .CP(n2114), .Q(n2075) );
  CFD1QX4 clk_r_REG277_S1 ( .D(n572), .CP(n2114), .Q(net171595) );
  CFD1QX2 clk_r_REG275_S1 ( .D(n478), .CP(n2114), .Q(n2068) );
  CFD1QX2 clk_r_REG205_S1 ( .D(n272), .CP(n2114), .Q(n2109) );
  CFD1QX2 clk_r_REG203_S1 ( .D(n277), .CP(n2114), .Q(n2107) );
  CFD1QX2 clk_r_REG189_S1 ( .D(n422), .CP(n2114), .Q(n2083) );
  CFD1QX2 clk_r_REG270_S1 ( .D(n520), .CP(n2114), .Q(n2059) );
  CFD1QX4 clk_r_REG178_S1 ( .D(n676), .CP(n2114), .Q(n2036) );
  CFD1QX2 clk_r_REG218_S1 ( .D(n521), .CP(n2114), .Q(n2096) );
  CFD1QX2 clk_r_REG193_S1 ( .D(n450), .CP(n2114), .Q(n2076) );
  CFD1QX2 clk_r_REG212_S1 ( .D(n524), .CP(n2114), .Q(n2057) );
  CFD1QX2 clk_r_REG222_S1 ( .D(n496), .CP(n2114), .Q(n2065) );
  CFD1QX1 clk_r_REG244_S1 ( .D(n369), .CP(n2114), .Q(n2101) );
  CFD1QX2 clk_r_REG182_S1 ( .D(n674), .CP(n2114), .Q(n2037) );
  CFD1QX2 clk_r_REG186_S1 ( .D(n445), .CP(n2114), .Q(n2081) );
  CFD1QX2 clk_r_REG263_S1 ( .D(n417), .CP(n2114), .Q(n2088) );
  CFD1QX2 clk_r_REG176_S1 ( .D(n688), .CP(n2114), .Q(n2034) );
  CFD1QX2 clk_r_REG269_S1 ( .D(n519), .CP(n2114), .Q(n2060) );
  CFD1QX2 clk_r_REG240_S1 ( .D(n424), .CP(n2114), .Q(n2082) );
  CFD1QX2 clk_r_REG259_S1 ( .D(n545), .CP(n2114), .Q(n2056) );
  CFD1QX2 clk_r_REG220_S1 ( .D(n500), .CP(n2114), .Q(n2061) );
  CFD1QX1 clk_r_REG227_S1 ( .D(n568), .CP(n2114), .Q(net171593) );
  CFD1QX2 clk_r_REG247_S1 ( .D(n475), .CP(n2114), .Q(n2070) );
  CFD1QX1 clk_r_REG223_S1 ( .D(n473), .CP(n2114), .Q(n2072) );
  CFD1QX1 clk_r_REG225_S1 ( .D(n585), .CP(n2114), .Q(net171600) );
  CFD1QX1 clk_r_REG253_S1 ( .D(n447), .CP(n2114), .Q(n2079) );
  CFD1QX2 clk_r_REG251_S1 ( .D(n588), .CP(n2114), .Q(n2053) );
  CFD1QX2 clk_r_REG215_S1 ( .D(n541), .CP(n2114), .Q(net171496) );
  CFD1QX2 clk_r_REG230_S1 ( .D(n584), .CP(n2114), .Q(net171599) );
  CFD1QX2 clk_r_REG246_S1 ( .D(n498), .CP(n2114), .Q(n2063) );
  CFA1X1 U486 ( .A(net171599), .B(n582), .CI(n601), .CO(n579), .S(n580) );
  CND2IX1 U601 ( .B(net33078), .A(a[31]), .Z(n1088) );
  CFD1QX2 clk_r_REG248_S1 ( .D(n476), .CP(n2114), .Q(n2069) );
  CFD1QX2 clk_r_REG190_S1 ( .D(n471), .CP(n2114), .Q(n2074) );
  CFD1QX2 clk_r_REG226_S1 ( .D(n586), .CP(n2114), .Q(n2054) );
  CEOX2 U1263 ( .A(a[0]), .B(net32098), .Z(n1421) );
  COND2X1 U1108 ( .A(n1548), .B(n1343), .C(n6), .D(n1342), .Z(n1056) );
  COND2X1 U1110 ( .A(n1548), .B(n1345), .C(n6), .D(n1344), .Z(n1058) );
  COND2X1 U605 ( .A(n112), .B(n1092), .C(n1091), .D(n110), .Z(n819) );
  CFD1QXL clk_r_REG228_S1 ( .D(n606), .CP(n2114), .Q(n2050) );
  CFD1QX2 clk_r_REG199_S1 ( .D(n286), .CP(n2114), .Q(n2104) );
  CFD1QX2 clk_r_REG209_S1 ( .D(n1813), .CP(n2114), .Q(n2113) );
  CFD1QX2 clk_r_REG200_S1 ( .D(n279), .CP(n2114), .Q(n2097) );
  CFD1QX2 clk_r_REG255_S1 ( .D(n419), .CP(n2114), .Q(n2086) );
  CFD1QX2 clk_r_REG238_S1 ( .D(n392), .CP(n2114), .Q(n2092) );
  CFD1QX2 clk_r_REG260_S1 ( .D(n546), .CP(n2114), .Q(net171589) );
  CFD1QX2 clk_r_REG229_S1 ( .D(n583), .CP(n2114), .Q(net171598) );
  CFD1QX2 clk_r_REG237_S1 ( .D(n391), .CP(n2114), .Q(n2093) );
  CFD1QX4 clk_r_REG278_S1 ( .D(n591), .CP(n2114), .Q(net171605) );
  CFD1QX1 clk_r_REG180_S1 ( .D(n658), .CP(n2114), .Q(n2040) );
  CFD1QX2 clk_r_REG214_S1 ( .D(n542), .CP(n2114), .Q(net171472) );
  CFD1QX2 clk_r_REG242_S1 ( .D(n390), .CP(n2114), .Q(n2094) );
  CFD1QX1 clk_r_REG185_S1 ( .D(n640), .CP(n2114), .Q(n2044) );
  CFD1QX2 clk_r_REG232_S1 ( .D(n628), .CP(n2114), .Q(n2046) );
  CFD1QX1 clk_r_REG194_S1 ( .D(n370), .CP(n2114), .Q(n2100) );
  CFD1QX2 clk_r_REG236_S1 ( .D(n608), .CP(n2114), .Q(n2049) );
  CFD1QX4 clk_r_REG177_S1 ( .D(n689), .CP(n2114), .Q(n2033) );
  CFD1QX2 clk_r_REG217_S1 ( .D(n522), .CP(n2114), .Q(n2102) );
  CFD1QX4 clk_r_REG252_S1 ( .D(n552), .CP(n2114), .Q(net171498) );
  CFD1QX2 clk_r_REG211_S1 ( .D(n523), .CP(n2114), .Q(n2058) );
  CFD1QX2 clk_r_REG264_S1 ( .D(n418), .CP(n2114), .Q(n2087) );
  CFD1QX2 clk_r_REG262_S1 ( .D(n482), .CP(n2114), .Q(n2067) );
  CFD1QX4 clk_r_REG276_S1 ( .D(n550), .CP(n2114), .Q(net171591) );
  CFD1QX4 clk_r_REG216_S1 ( .D(n547), .CP(n2114), .Q(n2055) );
  CFD1QX1 clk_r_REG191_S1 ( .D(n472), .CP(n2114), .Q(n2073) );
  CFD1QX2 clk_r_REG233_S1 ( .D(n603), .CP(n2114), .Q(n2052) );
  CFD1QX2 clk_r_REG234_S1 ( .D(n604), .CP(n2114), .Q(n2051) );
  CND2X4 U1267 ( .A(n1411), .B(n89), .Z(n91) );
  CNIVX1 U1268 ( .A(n852), .Z(n1666) );
  COND2X1 U1269 ( .A(n91), .B(n1129), .C(n89), .D(n1128), .Z(n852) );
  CENX2 U1270 ( .A(n127), .B(n215), .Z(product[23]) );
  COND1X2 U1271 ( .A(n216), .B(n222), .C(n1806), .Z(n215) );
  CENXL U1272 ( .A(n2151), .B(n2168), .Z(n1130) );
  CENXL U1273 ( .A(net33076), .B(n2168), .Z(n1132) );
  CENXL U1274 ( .A(net33422), .B(n2168), .Z(n1131) );
  CENXL U1275 ( .A(n2158), .B(n2168), .Z(n1123) );
  CENX1 U1276 ( .A(n2153), .B(n2168), .Z(n1128) );
  CND2X1 U1277 ( .A(n2118), .B(n1547), .Z(n1939) );
  CIVXL U1278 ( .A(n2107), .Z(n275) );
  CIVX1 U1279 ( .A(net180562), .Z(n1433) );
  CIVX1 U1280 ( .A(n1433), .Z(net182741) );
  CEOX1 U1281 ( .A(n887), .B(n857), .Z(n1543) );
  CEOX2 U1282 ( .A(n1543), .B(n821), .Z(n375) );
  COR2XL U1283 ( .A(n1095), .B(n107), .Z(n1544) );
  COR2XL U1284 ( .A(n1094), .B(n1812), .Z(n1545) );
  CND2X2 U1285 ( .A(n1544), .B(n1545), .Z(n821) );
  CENXL U1286 ( .A(n2153), .B(net182741), .Z(n1095) );
  CNIVX4 U1287 ( .A(n63), .Z(n2165) );
  COR2XL U1288 ( .A(n1096), .B(n107), .Z(n1877) );
  CIVX1 U1289 ( .A(n837), .Z(n1546) );
  CIVX2 U1290 ( .A(n1546), .Z(n1547) );
  CND2X1 U1291 ( .A(n1993), .B(n1994), .Z(product[21]) );
  CND2XL U1292 ( .A(n1407), .B(net184424), .Z(n1574) );
  CNIVX3 U1293 ( .A(n9), .Z(n1548) );
  CIVX1 U1294 ( .A(n882), .Z(n1549) );
  CIVX2 U1295 ( .A(n1549), .Z(n1550) );
  CEOXL U1296 ( .A(n1625), .B(n610), .Z(n604) );
  CIVX8 U1297 ( .A(n2182), .Z(n2178) );
  COND1X2 U1298 ( .A(n317), .B(n315), .C(n316), .Z(n314) );
  CANR1X2 U1299 ( .A(n322), .B(n2021), .C(n319), .Z(n317) );
  COND1X2 U1300 ( .A(n307), .B(n309), .C(n308), .Z(n306) );
  CANR1X2 U1301 ( .A(n314), .B(n2022), .C(n311), .Z(n309) );
  CEO3XL U1302 ( .A(n629), .B(n612), .C(n614), .Z(n606) );
  CIVX1 U1303 ( .A(n946), .Z(n1551) );
  CIVX1 U1304 ( .A(n1551), .Z(n1552) );
  CEO3XL U1305 ( .A(n732), .B(n730), .C(n741), .Z(n1553) );
  CND2IXL U1306 ( .B(net33078), .A(n2204), .Z(n1205) );
  COND2X1 U1307 ( .A(n61), .B(n1203), .C(n58), .D(n1202), .Z(n922) );
  CAN2X1 U1308 ( .A(n342), .B(n1806), .Z(net178962) );
  CIVDX1 U1309 ( .A(n217), .Z0(n1807), .Z1(n1806) );
  CENX2 U1310 ( .A(n1554), .B(n831), .Z(n480) );
  CENX1 U1311 ( .A(n951), .B(n975), .Z(n1554) );
  CFA1XL U1312 ( .A(n861), .B(n929), .CI(n875), .CO(n483), .S(n484) );
  CFA1XL U1313 ( .A(n904), .B(n922), .CI(n942), .CO(n725), .S(n726) );
  CIVXL U1314 ( .A(n719), .Z(n1847) );
  CFA1XL U1315 ( .A(n938), .B(n1038), .CI(n1010), .CO(n665), .S(n666) );
  CND2XL U1316 ( .A(n1958), .B(n1957), .Z(n1555) );
  CAOR1X1 U1317 ( .A(n2020), .B(n1968), .C(n154), .Z(n1556) );
  CND2XL U1318 ( .A(n1958), .B(n1957), .Z(n1968) );
  COR2X1 U1319 ( .A(n100), .B(n1104), .Z(n1948) );
  CND2X1 U1320 ( .A(n1644), .B(n1816), .Z(n53) );
  CND2IX2 U1321 ( .B(n1699), .A(n1973), .Z(n1974) );
  CNR2XL U1322 ( .A(n1986), .B(n167), .Z(n1557) );
  CNR2XL U1323 ( .A(n1986), .B(n167), .Z(n1558) );
  CND2XL U1324 ( .A(n953), .B(n802), .Z(n1559) );
  COND2XL U1325 ( .A(n2117), .B(n1224), .C(n1223), .D(n1815), .Z(n942) );
  CENXL U1326 ( .A(n1560), .B(n430), .Z(n418) );
  CENX1 U1327 ( .A(n428), .B(n426), .Z(n1560) );
  CND2IX2 U1328 ( .B(n953), .A(n1656), .Z(n1657) );
  CEO3XL U1329 ( .A(n466), .B(n464), .C(n489), .Z(n1561) );
  COR2X1 U1330 ( .A(n58), .B(n1201), .Z(n1884) );
  CENXL U1331 ( .A(n2152), .B(n2203), .Z(n1201) );
  CIVX1 U1332 ( .A(n194), .Z(n192) );
  CIVXL U1333 ( .A(n469), .Z(n1562) );
  CIVX1 U1334 ( .A(n1562), .Z(n1563) );
  CANR1X1 U1335 ( .A(n2020), .B(n1555), .C(n154), .Z(n1564) );
  CENX1 U1336 ( .A(n1783), .B(n1782), .Z(n1781) );
  CND2X1 U1337 ( .A(n1878), .B(n1877), .Z(n1565) );
  CND2X1 U1338 ( .A(n1878), .B(n1877), .Z(n822) );
  COR2XL U1339 ( .A(n1814), .B(n1105), .Z(n1844) );
  CEOX1 U1340 ( .A(n1632), .B(n921), .Z(n712) );
  CNR2IX1 U1341 ( .B(net33078), .A(n105), .Z(n826) );
  CENXL U1342 ( .A(n2152), .B(n1835), .Z(n1105) );
  CND2X2 U1343 ( .A(n1409), .B(n100), .Z(n102) );
  CIVX3 U1344 ( .A(net184082), .Z(net183987) );
  CIVXL U1345 ( .A(net184082), .Z(net183988) );
  CND2X2 U1346 ( .A(n1575), .B(n1948), .Z(n830) );
  CND2XL U1347 ( .A(n824), .B(n1745), .Z(n1568) );
  CND2X2 U1348 ( .A(n1566), .B(n1567), .Z(n1569) );
  CND2X2 U1349 ( .A(n1568), .B(n1569), .Z(n454) );
  CIVX1 U1350 ( .A(n824), .Z(n1566) );
  CIVX2 U1351 ( .A(n1745), .Z(n1567) );
  CIVX1 U1352 ( .A(n404), .Z(n1749) );
  CENX1 U1353 ( .A(net33076), .B(n1857), .Z(n1183) );
  COND1X1 U1354 ( .A(n184), .B(n178), .C(n179), .Z(n173) );
  COND2X1 U1355 ( .A(n1932), .B(n1182), .C(n66), .D(n1181), .Z(n902) );
  CENX4 U1356 ( .A(n278), .B(n137), .Z(product[13]) );
  CND2X4 U1357 ( .A(n1991), .B(n1990), .Z(product[29]) );
  COR2XL U1358 ( .A(n1097), .B(n107), .Z(n1616) );
  CND2IX1 U1359 ( .B(n2026), .A(n66), .Z(n1570) );
  CENX2 U1360 ( .A(net178513), .B(n514), .Z(n512) );
  CND2X2 U1361 ( .A(n1760), .B(n1759), .Z(n514) );
  CANR1X1 U1362 ( .A(net179842), .B(n1805), .C(n192), .Z(n190) );
  CND2X2 U1363 ( .A(n740), .B(n749), .Z(n283) );
  CND2X1 U1364 ( .A(n1974), .B(n1975), .Z(n1571) );
  CND2X2 U1365 ( .A(n1974), .B(n1975), .Z(n1409) );
  CEOX4 U1366 ( .A(n1654), .B(a[12]), .Z(n58) );
  CIVX1 U1367 ( .A(n920), .Z(n1572) );
  CIVX2 U1368 ( .A(n1572), .Z(n1573) );
  CND2X1 U1369 ( .A(n953), .B(n802), .Z(n1898) );
  CND2IX1 U1370 ( .B(n2026), .A(n66), .Z(n69) );
  CND2X2 U1371 ( .A(n431), .B(n998), .Z(n1680) );
  CND2XL U1372 ( .A(n1407), .B(net184424), .Z(net179858) );
  COR2X1 U1373 ( .A(n1105), .B(n102), .Z(n1575) );
  CIVXL U1374 ( .A(n1748), .Z(n1576) );
  CIVX2 U1375 ( .A(n406), .Z(n1748) );
  CIVX2 U1376 ( .A(n48), .Z(n1654) );
  CAN2X1 U1377 ( .A(n2104), .B(n2113), .Z(n1577) );
  CND2IX2 U1378 ( .B(n2105), .A(n1577), .Z(n1751) );
  CND2IX4 U1379 ( .B(n2113), .A(n139), .Z(n1752) );
  CND3X1 U1380 ( .A(n1940), .B(n1938), .C(n1939), .Z(n431) );
  CND3XL U1381 ( .A(n1938), .B(n1940), .C(n1939), .Z(n1578) );
  CND2XL U1382 ( .A(n1582), .B(n426), .Z(n1579) );
  CND2XL U1383 ( .A(n1582), .B(n428), .Z(n1580) );
  CND2XL U1384 ( .A(n426), .B(n428), .Z(n1581) );
  CND3XL U1385 ( .A(n1579), .B(n1580), .C(n1581), .Z(n417) );
  CENXL U1386 ( .A(n1618), .B(n823), .Z(n1582) );
  CND2X2 U1387 ( .A(n1621), .B(n1622), .Z(n428) );
  CENXL U1388 ( .A(n1618), .B(n823), .Z(n430) );
  CND2X1 U1389 ( .A(n1616), .B(n1617), .Z(n823) );
  CND2X1 U1390 ( .A(n800), .B(n2118), .Z(n1938) );
  CENX1 U1391 ( .A(net33422), .B(net180562), .Z(n1098) );
  CNIVX3 U1392 ( .A(n63), .Z(n1856) );
  CHA1X2 U1393 ( .A(n807), .B(n963), .CO(n713), .S(n714) );
  CENX1 U1394 ( .A(n2157), .B(n1933), .Z(n1111) );
  CND2XL U1395 ( .A(net182672), .B(net183987), .Z(n1624) );
  CND3X2 U1396 ( .A(net179429), .B(net179428), .C(net179427), .Z(n543) );
  CND2X1 U1397 ( .A(net171591), .B(net171592), .Z(net179427) );
  CND2X1 U1398 ( .A(net171498), .B(net171592), .Z(net179429) );
  CENX1 U1399 ( .A(a[28]), .B(n1623), .Z(n110) );
  CENX1 U1400 ( .A(n1858), .B(n400), .Z(n392) );
  CND2XL U1401 ( .A(n819), .B(n1057), .Z(net179942) );
  CND2XL U1402 ( .A(n819), .B(n973), .Z(net179941) );
  CNR2X2 U1403 ( .A(n1961), .B(n2035), .Z(n251) );
  CND2X1 U1404 ( .A(net171591), .B(net171498), .Z(net179428) );
  CND2X1 U1405 ( .A(n1775), .B(n1779), .Z(n1759) );
  CENX2 U1406 ( .A(net171498), .B(net171591), .Z(n1782) );
  CND3X2 U1407 ( .A(n1776), .B(n1778), .C(n1777), .Z(n1775) );
  CND2X1 U1408 ( .A(n1801), .B(n1795), .Z(n1776) );
  CND2X1 U1409 ( .A(n1801), .B(net171589), .Z(n1778) );
  CND2X1 U1410 ( .A(n1780), .B(n1792), .Z(n1760) );
  CND2X1 U1411 ( .A(net171600), .B(net171602), .Z(n1800) );
  CENX1 U1412 ( .A(net171600), .B(net171593), .Z(n1790) );
  CNR2IX1 U1413 ( .B(n1779), .A(n1780), .Z(n1763) );
  CND3XL U1414 ( .A(n1796), .B(n1803), .C(n1802), .Z(n1761) );
  CND2XL U1415 ( .A(n1786), .B(n1787), .Z(n1802) );
  CND2X1 U1416 ( .A(net33776), .B(n1794), .Z(n1789) );
  CND2X1 U1417 ( .A(n1793), .B(n1797), .Z(n1794) );
  CND2XL U1418 ( .A(n581), .B(n1583), .Z(net179824) );
  CND2XL U1419 ( .A(n560), .B(n1583), .Z(net179825) );
  CND2XL U1420 ( .A(n581), .B(n560), .Z(n1949) );
  CND2X1 U1421 ( .A(n2069), .B(n2071), .Z(n1642) );
  CND2X1 U1422 ( .A(n2064), .B(n2071), .Z(n1643) );
  CANR1X1 U1423 ( .A(net178512), .B(n232), .C(n227), .Z(n225) );
  CENX1 U1424 ( .A(n516), .B(n1761), .Z(net178513) );
  CND2X1 U1425 ( .A(n136), .B(n1638), .Z(n1639) );
  CND2X1 U1426 ( .A(n164), .B(n2016), .Z(n1990) );
  CENX1 U1427 ( .A(n253), .B(n133), .Z(product[17]) );
  COND1X1 U1428 ( .A(n254), .B(n260), .C(n255), .Z(n253) );
  CIVX2 U1429 ( .A(n12), .Z(n2175) );
  CIVX4 U1430 ( .A(n1654), .Z(n2200) );
  CEOX1 U1431 ( .A(n1071), .B(n941), .Z(n1632) );
  CND2X1 U1432 ( .A(n1735), .B(a[31]), .Z(n1733) );
  CND2X1 U1433 ( .A(n801), .B(n839), .Z(n1704) );
  CND2IX2 U1434 ( .B(n2012), .A(n42), .Z(n44) );
  CNR2X1 U1435 ( .A(n1608), .B(n749), .Z(n282) );
  CENX1 U1436 ( .A(n453), .B(n451), .Z(n1655) );
  CIVX2 U1437 ( .A(n549), .Z(n1895) );
  CEOX2 U1438 ( .A(n1790), .B(n1771), .Z(n1583) );
  CNIVX1 U1439 ( .A(n910), .Z(n1584) );
  CNIVX1 U1440 ( .A(n1932), .Z(n1585) );
  CNIVX1 U1441 ( .A(n1697), .Z(n1586) );
  CNIVX1 U1442 ( .A(a[20]), .Z(n1587) );
  CIVX2 U1443 ( .A(n2168), .Z(n1436) );
  CEO3X1 U1444 ( .A(net171472), .B(n1786), .C(n1787), .Z(n1588) );
  CIVX1 U1445 ( .A(n30), .Z(n2189) );
  CIVX2 U1446 ( .A(n2189), .Z(n2183) );
  CAN3X1 U1447 ( .A(net179824), .B(net179825), .C(n1949), .Z(n1589) );
  CIVDXL U1448 ( .A(n183), .Z0(n1590), .Z1(n1591) );
  COR2X1 U1449 ( .A(n379), .B(n364), .Z(n1592) );
  COR2XL U1450 ( .A(n1085), .B(n814), .Z(n1593) );
  CANR1X2 U1451 ( .A(n2017), .B(n306), .C(n303), .Z(n301) );
  CIVX2 U1452 ( .A(n301), .Z(n300) );
  CNIVX2 U1453 ( .A(n79), .Z(n2167) );
  CENX1 U1454 ( .A(n423), .B(n398), .Z(n1597) );
  CENXL U1455 ( .A(n1597), .B(n402), .Z(n390) );
  CENX1 U1456 ( .A(n1594), .B(n662), .Z(n658) );
  CENX2 U1457 ( .A(n664), .B(n675), .Z(n1594) );
  CIVXL U1458 ( .A(n66), .Z(n1595) );
  CIVX1 U1459 ( .A(n1595), .Z(n1596) );
  CIVX4 U1460 ( .A(n2190), .Z(n2187) );
  CIVXL U1461 ( .A(n61), .Z(n1598) );
  CIVXL U1462 ( .A(n1598), .Z(n1599) );
  CNR2X1 U1463 ( .A(net171597), .B(net171605), .Z(n1767) );
  CND2X1 U1464 ( .A(net171605), .B(net171597), .Z(n1798) );
  CEOXL U1465 ( .A(n1864), .B(n616), .Z(n608) );
  CND2X4 U1466 ( .A(n1412), .B(n82), .Z(n84) );
  CENX1 U1467 ( .A(net33422), .B(n2138), .Z(n1146) );
  COND2XL U1468 ( .A(n44), .B(n1237), .C(n1236), .D(n42), .Z(n954) );
  COND2XL U1469 ( .A(n44), .B(n1238), .C(n1237), .D(n42), .Z(n955) );
  COND2XL U1470 ( .A(n44), .B(n1241), .C(n1240), .D(n42), .Z(n958) );
  COND2XL U1471 ( .A(n44), .B(n1239), .C(n1238), .D(n42), .Z(n956) );
  COND2XL U1472 ( .A(n44), .B(n1243), .C(n1242), .D(n42), .Z(n960) );
  COND2XL U1473 ( .A(n44), .B(n1245), .C(n1244), .D(n42), .Z(n962) );
  CNR2IXL U1474 ( .B(net33078), .A(n42), .Z(n970) );
  COND2XL U1475 ( .A(n44), .B(n1249), .C(n1248), .D(n42), .Z(n966) );
  COND2XL U1476 ( .A(n44), .B(n1250), .C(n1249), .D(n42), .Z(n967) );
  CENXL U1477 ( .A(n429), .B(n1600), .Z(n394) );
  CENX2 U1478 ( .A(n427), .B(n425), .Z(n1600) );
  CND3X2 U1479 ( .A(n1907), .B(n1908), .C(n1909), .Z(n427) );
  CIVX2 U1480 ( .A(n2166), .Z(n1935) );
  CENX2 U1481 ( .A(a[8]), .B(n2195), .Z(n2012) );
  CIVX3 U1482 ( .A(n2199), .Z(n2195) );
  CIVX1 U1483 ( .A(n186), .Z(net179617) );
  CEO3X1 U1484 ( .A(n948), .B(n888), .C(n1565), .Z(n400) );
  CNR2X2 U1485 ( .A(n1437), .B(n84), .Z(n1744) );
  COND2X1 U1486 ( .A(n1586), .B(n1156), .C(n74), .D(n1155), .Z(n877) );
  CFA1X1 U1487 ( .A(n931), .B(n851), .CI(n877), .CO(n531), .S(n532) );
  CEOX1 U1488 ( .A(n1739), .B(n652), .Z(n644) );
  CND2XL U1489 ( .A(n652), .B(n665), .Z(n1741) );
  CND2XL U1490 ( .A(n652), .B(n650), .Z(n1740) );
  CENX1 U1491 ( .A(n1601), .B(n602), .Z(n600) );
  CENX2 U1492 ( .A(n2051), .B(n621), .Z(n1601) );
  CEO3X1 U1493 ( .A(net171598), .B(n566), .C(n1756), .Z(n1791) );
  CIVX2 U1494 ( .A(a[24]), .Z(n1699) );
  CND2X2 U1495 ( .A(n1571), .B(n100), .Z(n1747) );
  CIVX2 U1496 ( .A(n55), .Z(n2205) );
  CENXL U1497 ( .A(net180562), .B(n2151), .Z(n1097) );
  COND2XL U1498 ( .A(n1586), .B(n1155), .C(n74), .D(n1154), .Z(n1602) );
  CENXL U1499 ( .A(n1603), .B(n832), .Z(n506) );
  CENX1 U1500 ( .A(n952), .B(n876), .Z(n1603) );
  CND3X2 U1501 ( .A(net33755), .B(n2150), .C(net33757), .Z(n511) );
  COND1X1 U1502 ( .A(n1762), .B(n1763), .C(n1761), .Z(net33757) );
  CENXL U1503 ( .A(n1604), .B(n295), .Z(product[10]) );
  CAN2X1 U1504 ( .A(n2018), .B(n294), .Z(n1604) );
  CND3XL U1505 ( .A(net33752), .B(n2149), .C(net33754), .Z(n1605) );
  CIVX2 U1506 ( .A(n186), .Z(n185) );
  CNIVX2 U1507 ( .A(n848), .Z(n1606) );
  CAOR1XL U1508 ( .A(n261), .B(n242), .C(n243), .Z(n1661) );
  CND2X1 U1509 ( .A(n1698), .B(n1699), .Z(n1701) );
  COND2X1 U1510 ( .A(n1133), .B(n89), .C(n1436), .D(n91), .Z(n1607) );
  COND2XL U1511 ( .A(n1133), .B(n89), .C(n1436), .D(n91), .Z(n804) );
  COND2XL U1512 ( .A(n18), .B(n1334), .C(n1333), .D(n15), .Z(n1048) );
  CENX1 U1513 ( .A(n2171), .B(n2155), .Z(n1333) );
  CEO3XL U1514 ( .A(n751), .B(n744), .C(n742), .Z(n1608) );
  CND2X1 U1515 ( .A(net178512), .B(n229), .Z(n129) );
  COND1XL U1516 ( .A(n184), .B(n1611), .C(n179), .Z(n1609) );
  COND1XL U1517 ( .A(n184), .B(n1611), .C(n179), .Z(n1682) );
  CND3X2 U1518 ( .A(n1825), .B(n1826), .C(n1827), .Z(n709) );
  COND1X1 U1519 ( .A(n205), .B(n222), .C(net178660), .Z(n2004) );
  CANR1X2 U1520 ( .A(n351), .B(n278), .C(n275), .Z(n273) );
  CIVX3 U1521 ( .A(n2097), .Z(n278) );
  CND2X2 U1522 ( .A(n1556), .B(n119), .Z(n2014) );
  COND2X1 U1523 ( .A(n36), .B(n1274), .C(n1273), .D(net178746), .Z(n990) );
  CFA1X1 U1524 ( .A(n990), .B(n1074), .CI(n1044), .CO(n745), .S(n746) );
  CENXL U1525 ( .A(n1845), .B(n460), .Z(n448) );
  CND2XL U1526 ( .A(n833), .B(n1003), .Z(n1674) );
  CND2XL U1527 ( .A(n833), .B(n1031), .Z(n1675) );
  CEOX2 U1528 ( .A(n1673), .B(n833), .Z(n526) );
  CND3X1 U1529 ( .A(n1674), .B(n1675), .C(n1676), .Z(n525) );
  COND2XL U1530 ( .A(n1585), .B(n1177), .C(n66), .D(n1176), .Z(n897) );
  CNIVX4 U1531 ( .A(n86), .Z(n2168) );
  CNR2XL U1532 ( .A(n282), .B(n285), .Z(n280) );
  CNR2X1 U1533 ( .A(n487), .B(n1561), .Z(n1610) );
  CNR2XL U1534 ( .A(n462), .B(n487), .Z(n1611) );
  CNR2X1 U1535 ( .A(n1561), .B(n487), .Z(n178) );
  CND2X2 U1536 ( .A(n1919), .B(n1920), .Z(product[18]) );
  CNR2IX1 U1537 ( .B(net33078), .A(n110), .Z(n820) );
  CIVXL U1538 ( .A(n223), .Z(n1612) );
  CIVXL U1539 ( .A(n490), .Z(n1613) );
  CIVX1 U1540 ( .A(n1613), .Z(n1614) );
  CND3X2 U1541 ( .A(n1679), .B(n1680), .C(n1681), .Z(n395) );
  CND2XL U1542 ( .A(n1576), .B(n404), .Z(n1615) );
  CENX1 U1543 ( .A(net184434), .B(n819), .Z(n426) );
  CENX1 U1544 ( .A(n1057), .B(n973), .Z(net184434) );
  CENXL U1545 ( .A(n907), .B(n859), .Z(n1618) );
  CND2XL U1546 ( .A(n1619), .B(n829), .Z(n1622) );
  CIVXL U1547 ( .A(net180068), .Z(n1619) );
  CND2X1 U1548 ( .A(net180068), .B(n1620), .Z(n1621) );
  CIVXL U1549 ( .A(n829), .Z(n1620) );
  CENXL U1550 ( .A(net33076), .B(net183987), .Z(n1092) );
  CIVX2 U1551 ( .A(n109), .Z(net184082) );
  CNIVX2 U1552 ( .A(n116), .Z(net33076) );
  COND2XL U1553 ( .A(n1548), .B(n1344), .C(n6), .D(n1343), .Z(n1057) );
  CND2X1 U1554 ( .A(n973), .B(n1057), .Z(net179943) );
  CIVX4 U1555 ( .A(a[0]), .Z(n6) );
  COND2XL U1556 ( .A(n36), .B(n1257), .C(n1256), .D(net178746), .Z(n973) );
  CND2XL U1557 ( .A(n823), .B(n907), .Z(net180365) );
  CND2XL U1558 ( .A(n823), .B(n859), .Z(net180364) );
  COR2XL U1559 ( .A(net181698), .B(n1096), .Z(n1617) );
  COND2XL U1560 ( .A(n1599), .B(n1188), .C(n1187), .D(net180674), .Z(n907) );
  CND2XL U1561 ( .A(n859), .B(n907), .Z(net180366) );
  CND2X1 U1562 ( .A(n1407), .B(net184424), .Z(n112) );
  COR2XL U1563 ( .A(n1091), .B(n112), .Z(net180011) );
  CND2X1 U1564 ( .A(n1624), .B(net182674), .Z(n1407) );
  CIVX2 U1565 ( .A(a[28]), .Z(net182672) );
  CND2XL U1566 ( .A(net182673), .B(a[28]), .Z(net182674) );
  CIVXL U1567 ( .A(net183988), .Z(net182673) );
  CNIVX4 U1568 ( .A(n104), .Z(n1623) );
  CENX2 U1569 ( .A(a[28]), .B(n1623), .Z(net184424) );
  CNIVX4 U1570 ( .A(n104), .Z(net180562) );
  CNIVX4 U1571 ( .A(n116), .Z(net33078) );
  COND2XL U1572 ( .A(n36), .B(n1258), .C(n1257), .D(net178746), .Z(n974) );
  COND2XL U1573 ( .A(n36), .B(n1256), .C(n1255), .D(net178746), .Z(n972) );
  CENXL U1574 ( .A(net33422), .B(net183987), .Z(n1091) );
  CNIVX4 U1575 ( .A(n1404), .Z(net33422) );
  CEOX1 U1576 ( .A(n1653), .B(n818), .Z(n402) );
  COND2X1 U1577 ( .A(n1116), .B(n97), .C(n95), .D(n1115), .Z(n840) );
  CEO3X2 U1578 ( .A(n1007), .B(n635), .C(n618), .Z(n610) );
  CEOX2 U1579 ( .A(n627), .B(n625), .Z(n1625) );
  CND2XL U1580 ( .A(n1007), .B(n635), .Z(n1626) );
  CND2X1 U1581 ( .A(n1007), .B(n618), .Z(n1627) );
  CND2XL U1582 ( .A(n635), .B(n618), .Z(n1628) );
  CND3X1 U1583 ( .A(n1626), .B(n1627), .C(n1628), .Z(n609) );
  CND2XL U1584 ( .A(n627), .B(n625), .Z(n1629) );
  CND2XL U1585 ( .A(n627), .B(n610), .Z(n1630) );
  CND2XL U1586 ( .A(n625), .B(n610), .Z(n1631) );
  CND3XL U1587 ( .A(n1629), .B(n1630), .C(n1631), .Z(n603) );
  CENXL U1588 ( .A(n2195), .B(n1388), .Z(n1235) );
  CENXL U1589 ( .A(net33076), .B(n2195), .Z(n1252) );
  CENXL U1590 ( .A(net33422), .B(n2195), .Z(n1251) );
  CND2X1 U1591 ( .A(n921), .B(n941), .Z(n1633) );
  CND2X1 U1592 ( .A(n921), .B(n1071), .Z(n1634) );
  CND2XL U1593 ( .A(n941), .B(n1071), .Z(n1635) );
  CND3X2 U1594 ( .A(n1633), .B(n1634), .C(n1635), .Z(n711) );
  COND1X1 U1595 ( .A(n167), .B(n175), .C(n170), .Z(n1636) );
  CNR2X2 U1596 ( .A(n436), .B(n461), .Z(n167) );
  COND1X1 U1597 ( .A(n167), .B(n175), .C(n170), .Z(n166) );
  CND2X1 U1598 ( .A(n1564), .B(n2013), .Z(n2015) );
  CANR1XL U1599 ( .A(n1682), .B(n1557), .C(n161), .Z(n159) );
  CEOX1 U1600 ( .A(n1953), .B(n1563), .Z(n440) );
  CND2X1 U1601 ( .A(n1637), .B(n273), .Z(n1640) );
  CND2X2 U1602 ( .A(n1639), .B(n1640), .Z(product[14]) );
  CIVX1 U1603 ( .A(n136), .Z(n1637) );
  CIVX2 U1604 ( .A(n273), .Z(n1638) );
  CEO3X1 U1605 ( .A(n2069), .B(n2071), .C(n2064), .Z(n468) );
  CND2X1 U1606 ( .A(n2069), .B(n2064), .Z(n1641) );
  CND3X2 U1607 ( .A(n1641), .B(n1642), .C(n1643), .Z(n467) );
  CEOX2 U1608 ( .A(n2080), .B(n467), .Z(n1953) );
  CENXL U1609 ( .A(a[10]), .B(n1654), .Z(n1644) );
  CEO3X2 U1610 ( .A(n681), .B(n670), .C(n668), .Z(n662) );
  CND2XL U1611 ( .A(n681), .B(n670), .Z(n1645) );
  CND2X1 U1612 ( .A(n681), .B(n668), .Z(n1646) );
  CND2X1 U1613 ( .A(n670), .B(n668), .Z(n1647) );
  CND3X1 U1614 ( .A(n1645), .B(n1646), .C(n1647), .Z(n661) );
  CND2XL U1615 ( .A(n664), .B(n675), .Z(n1648) );
  CND2XL U1616 ( .A(n664), .B(n662), .Z(n1649) );
  CND2XL U1617 ( .A(n675), .B(n662), .Z(n1650) );
  CND3XL U1618 ( .A(n1648), .B(n1649), .C(n1650), .Z(n657) );
  CEOX2 U1619 ( .A(n456), .B(n1944), .Z(n446) );
  COR2X1 U1620 ( .A(n97), .B(n1111), .Z(n1651) );
  COR2XL U1621 ( .A(n95), .B(n1110), .Z(n1652) );
  CND2X2 U1622 ( .A(n1651), .B(n1652), .Z(n835) );
  CEO3X1 U1623 ( .A(n905), .B(n835), .C(n799), .Z(n377) );
  CIVXL U1624 ( .A(n1760), .Z(n1762) );
  CEOX1 U1625 ( .A(n906), .B(n858), .Z(n1653) );
  CND2X1 U1626 ( .A(net180011), .B(n1927), .Z(n818) );
  CND3X2 U1627 ( .A(net179941), .B(net179942), .C(net179943), .Z(n425) );
  CND2IX1 U1628 ( .B(n1662), .A(n1995), .Z(n1997) );
  CND2X1 U1629 ( .A(n903), .B(n1041), .Z(n1826) );
  CND2X1 U1630 ( .A(n903), .B(n987), .Z(n1825) );
  CND2X2 U1631 ( .A(n1981), .B(n1436), .Z(n1983) );
  CNR2IX2 U1632 ( .B(net33078), .A(n1729), .Z(n816) );
  CIVX8 U1633 ( .A(n21), .Z(n2182) );
  COND2X1 U1634 ( .A(n36), .B(n1278), .C(n1277), .D(net178746), .Z(n994) );
  COND2XL U1635 ( .A(n1585), .B(n1172), .C(n1596), .D(n1171), .Z(n892) );
  CNR2IX1 U1636 ( .B(net33078), .A(n66), .Z(n904) );
  CENXL U1637 ( .A(n432), .B(n1655), .Z(n420) );
  CND2X2 U1638 ( .A(n1997), .B(n1996), .Z(product[19]) );
  CHA1XL U1639 ( .A(n901), .B(n939), .CO(n685), .S(n686) );
  CND2X2 U1640 ( .A(n1898), .B(n1657), .Z(n1671) );
  CIVX2 U1641 ( .A(n802), .Z(n1656) );
  COND2X1 U1642 ( .A(n1118), .B(n97), .C(n95), .D(n1117), .Z(n842) );
  CND2XL U1643 ( .A(n93), .B(a[24]), .Z(n1659) );
  CND2X1 U1644 ( .A(n1658), .B(n1698), .Z(n1660) );
  CND2X2 U1645 ( .A(n1659), .B(n1660), .Z(n100) );
  CIVXL U1646 ( .A(a[24]), .Z(n1658) );
  CAOR1X2 U1647 ( .A(n261), .B(n242), .C(n243), .Z(n1662) );
  CENX2 U1648 ( .A(n1663), .B(n615), .Z(n590) );
  CENX1 U1649 ( .A(n613), .B(n617), .Z(n1663) );
  CHA1X1 U1650 ( .A(n867), .B(n897), .CO(n617), .S(n618) );
  COND2X1 U1651 ( .A(n84), .B(n1145), .C(n82), .D(n1144), .Z(n867) );
  CND2X1 U1652 ( .A(n1992), .B(n129), .Z(n1993) );
  CND2IX1 U1653 ( .B(n158), .A(net179617), .Z(n1958) );
  CIVX1 U1654 ( .A(n566), .Z(n1754) );
  CENX2 U1655 ( .A(n1804), .B(net171605), .Z(n566) );
  CENX1 U1656 ( .A(n2156), .B(n1933), .Z(n1112) );
  CEO3XL U1657 ( .A(n492), .B(n1605), .C(n1614), .Z(n1664) );
  CIVX4 U1658 ( .A(n2202), .Z(n2201) );
  CNIVX2 U1659 ( .A(n993), .Z(n1665) );
  COR2X1 U1660 ( .A(n1977), .B(n1976), .Z(n944) );
  CNR2X1 U1661 ( .A(n2117), .B(n1226), .Z(n1976) );
  CNIVX2 U1662 ( .A(n1049), .Z(n1667) );
  CENXL U1663 ( .A(n2151), .B(n2201), .Z(n1668) );
  CND2XL U1664 ( .A(n1758), .B(n1588), .Z(net33775) );
  CIVX1 U1665 ( .A(n1758), .Z(n1793) );
  CNR2X1 U1666 ( .A(n244), .B(n247), .Z(n242) );
  COND2XL U1667 ( .A(n1183), .B(n1932), .C(n66), .D(n1182), .Z(n1669) );
  CENX1 U1668 ( .A(net33422), .B(n1857), .Z(n1182) );
  COND2XL U1669 ( .A(n97), .B(n1115), .C(n95), .D(n1114), .Z(n839) );
  CNR2IX2 U1670 ( .B(net33078), .A(n95), .Z(n844) );
  CANR1XL U1671 ( .A(n1609), .B(n1557), .C(n161), .Z(n1670) );
  COND1X1 U1672 ( .A(n170), .B(n1986), .C(n163), .Z(n161) );
  CENX2 U1673 ( .A(n1899), .B(n1671), .Z(n530) );
  CNIVX4 U1674 ( .A(n71), .Z(n1672) );
  CND2XL U1675 ( .A(n654), .B(n669), .Z(n1723) );
  CND3X1 U1676 ( .A(n1896), .B(n1897), .C(n1559), .Z(n529) );
  CND3X2 U1677 ( .A(n2143), .B(n2144), .C(n2145), .Z(n625) );
  CEOX1 U1678 ( .A(n1031), .B(n1003), .Z(n1673) );
  CND2X1 U1679 ( .A(n1003), .B(n1031), .Z(n1676) );
  COND2XL U1680 ( .A(n27), .B(n1288), .C(n1287), .D(n24), .Z(n1003) );
  COND2XL U1681 ( .A(n18), .B(n1317), .C(n1316), .D(n15), .Z(n1031) );
  CND2XL U1682 ( .A(n1958), .B(n1670), .Z(n1677) );
  CEOX1 U1683 ( .A(n998), .B(n433), .Z(n1678) );
  CEOXL U1684 ( .A(n431), .B(n1678), .Z(n396) );
  CND2X1 U1685 ( .A(n1578), .B(n433), .Z(n1679) );
  CND2X1 U1686 ( .A(n433), .B(n998), .Z(n1681) );
  CND2X1 U1687 ( .A(n347), .B(n348), .Z(n247) );
  CEOX2 U1688 ( .A(n706), .B(n717), .Z(n1683) );
  CEOX2 U1689 ( .A(n1683), .B(n704), .Z(n702) );
  CND2XL U1690 ( .A(n704), .B(n717), .Z(n1684) );
  CND2XL U1691 ( .A(n704), .B(n706), .Z(n1685) );
  CND2XL U1692 ( .A(n717), .B(n706), .Z(n1686) );
  CND3XL U1693 ( .A(n1684), .B(n1685), .C(n1686), .Z(n701) );
  CND2X1 U1694 ( .A(n1900), .B(n1688), .Z(n1689) );
  CND2X2 U1695 ( .A(n1687), .B(n708), .Z(n1690) );
  CND2X2 U1696 ( .A(n1689), .B(n1690), .Z(n704) );
  CIVX2 U1697 ( .A(n1900), .Z(n1687) );
  CIVXL U1698 ( .A(n708), .Z(n1688) );
  CND2X1 U1699 ( .A(n2203), .B(a[14]), .Z(n1693) );
  CND2X2 U1700 ( .A(n1691), .B(n1692), .Z(n1694) );
  CND2X4 U1701 ( .A(n1693), .B(n1694), .Z(n66) );
  CIVX2 U1702 ( .A(n2203), .Z(n1691) );
  CIVX2 U1703 ( .A(a[14]), .Z(n1692) );
  CND2XL U1704 ( .A(n702), .B(n715), .Z(n267) );
  CENX1 U1705 ( .A(net33422), .B(n1835), .Z(n1737) );
  CENXL U1706 ( .A(n2151), .B(n2203), .Z(n1695) );
  CIVXL U1707 ( .A(n2205), .Z(n1696) );
  CIVX1 U1708 ( .A(n251), .Z(n347) );
  COND1X2 U1709 ( .A(n224), .B(n1808), .C(n225), .Z(n223) );
  CND2X2 U1710 ( .A(n2009), .B(n74), .Z(n1697) );
  CND2X2 U1711 ( .A(n1936), .B(n1937), .Z(n2009) );
  COR2X1 U1712 ( .A(n1812), .B(n1095), .Z(n1878) );
  COND2X1 U1713 ( .A(n91), .B(n1128), .C(n89), .D(n1127), .Z(n851) );
  CENX1 U1714 ( .A(net33422), .B(n2201), .Z(n1226) );
  CND2X2 U1715 ( .A(n2020), .B(n156), .Z(n120) );
  CND2XL U1716 ( .A(n93), .B(a[24]), .Z(n1700) );
  CND2X2 U1717 ( .A(n1700), .B(n1701), .Z(n1814) );
  CIVXL U1718 ( .A(n93), .Z(n1698) );
  CNR2IX2 U1719 ( .B(net33078), .A(n1814), .Z(n834) );
  CND2X1 U1720 ( .A(n160), .B(n172), .Z(n158) );
  CEO3XL U1721 ( .A(n909), .B(n801), .C(n839), .Z(n482) );
  CND2X1 U1722 ( .A(n909), .B(n801), .Z(n1702) );
  CND2X1 U1723 ( .A(n909), .B(n839), .Z(n1703) );
  CND3X2 U1724 ( .A(n1702), .B(n1703), .C(n1704), .Z(n481) );
  CEOX1 U1725 ( .A(n485), .B(n483), .Z(n1705) );
  CEOX2 U1726 ( .A(n1705), .B(n481), .Z(n450) );
  CND2XL U1727 ( .A(n485), .B(n483), .Z(n1706) );
  CND2X1 U1728 ( .A(n485), .B(n481), .Z(n1707) );
  CND2X1 U1729 ( .A(n483), .B(n481), .Z(n1708) );
  CND3X1 U1730 ( .A(n1706), .B(n1707), .C(n1708), .Z(n449) );
  CFA1X1 U1731 ( .A(n937), .B(n1067), .CI(n1009), .CO(n649), .S(n650) );
  COND2X1 U1732 ( .A(n53), .B(n1219), .C(n1218), .D(n1816), .Z(n937) );
  CIVXL U1733 ( .A(n61), .Z(net184277) );
  CIVX1 U1734 ( .A(net184277), .Z(net184278) );
  CEOX1 U1735 ( .A(n518), .B(net171496), .Z(n1792) );
  CENX1 U1736 ( .A(n518), .B(net171496), .Z(n1779) );
  CEO3X1 U1737 ( .A(n844), .B(n854), .C(n866), .Z(n598) );
  CND2XL U1738 ( .A(n844), .B(n854), .Z(n1709) );
  CND2XL U1739 ( .A(n844), .B(n866), .Z(n1710) );
  CND2XL U1740 ( .A(n854), .B(n866), .Z(n1711) );
  CND3X1 U1741 ( .A(n1709), .B(n1710), .C(n1711), .Z(n597) );
  CEOXL U1742 ( .A(n593), .B(n595), .Z(n1712) );
  CEOXL U1743 ( .A(n1712), .B(n597), .Z(n568) );
  CND2XL U1744 ( .A(n593), .B(n595), .Z(n1713) );
  CND2XL U1745 ( .A(n593), .B(n597), .Z(n1714) );
  CND2XL U1746 ( .A(n595), .B(n597), .Z(n1715) );
  CND3X1 U1747 ( .A(n1713), .B(n1714), .C(n1715), .Z(n567) );
  CND2X1 U1748 ( .A(n800), .B(n1547), .Z(n1940) );
  CND2X1 U1749 ( .A(n710), .B(n1847), .Z(n1848) );
  CND2X1 U1750 ( .A(n710), .B(n708), .Z(n1905) );
  CIVX1 U1751 ( .A(net179546), .Z(net179547) );
  CNIVX4 U1752 ( .A(n99), .Z(n2169) );
  CIVX1 U1753 ( .A(n261), .Z(n260) );
  CND2X1 U1754 ( .A(n408), .B(n435), .Z(n163) );
  CND3X1 U1755 ( .A(n1910), .B(n1911), .C(n1912), .Z(n453) );
  CFA1X1 U1756 ( .A(n886), .B(n902), .CI(n1573), .CO(n699), .S(n700) );
  CNR2IX1 U1757 ( .B(net33078), .A(n74), .Z(n886) );
  CEO3X2 U1758 ( .A(n2049), .B(n2048), .C(n2050), .Z(n602) );
  CND2X1 U1759 ( .A(n2049), .B(n2048), .Z(n1716) );
  CND2X1 U1760 ( .A(n2049), .B(n2050), .Z(n1717) );
  CND2X1 U1761 ( .A(n2048), .B(n2050), .Z(n1718) );
  CND3X2 U1762 ( .A(n1716), .B(n1717), .C(n1718), .Z(n601) );
  CND2XL U1763 ( .A(n2051), .B(n621), .Z(n1719) );
  CND2XL U1764 ( .A(n2051), .B(n602), .Z(n1720) );
  CND2XL U1765 ( .A(n621), .B(n602), .Z(n1721) );
  CND3X1 U1766 ( .A(n1719), .B(n1720), .C(n1721), .Z(n599) );
  CEOX1 U1767 ( .A(n669), .B(n667), .Z(n1722) );
  CEOX1 U1768 ( .A(n1722), .B(n654), .Z(n646) );
  CND2X1 U1769 ( .A(n654), .B(n667), .Z(n1724) );
  CND2XL U1770 ( .A(n669), .B(n667), .Z(n1725) );
  CND3XL U1771 ( .A(n1723), .B(n1724), .C(n1725), .Z(n645) );
  CAOR1X1 U1772 ( .A(n165), .B(n185), .C(n166), .Z(n1726) );
  CNR2IX1 U1773 ( .B(n172), .A(n167), .Z(n165) );
  CEOX1 U1774 ( .A(n397), .B(n378), .Z(n1727) );
  CEOXL U1775 ( .A(n401), .B(n1727), .Z(n371) );
  CND3XL U1776 ( .A(n1921), .B(n1922), .C(n1923), .Z(n401) );
  COND2X2 U1777 ( .A(n1093), .B(net179547), .C(n1432), .D(n1574), .Z(n800) );
  COND1XL U1778 ( .A(n2110), .B(n2107), .C(n2109), .Z(n1728) );
  CIVX1 U1779 ( .A(n1662), .Z(n1808) );
  COND1X1 U1780 ( .A(n244), .B(n248), .C(n245), .Z(n243) );
  CENX1 U1781 ( .A(n569), .B(n567), .Z(n2008) );
  CENX1 U1782 ( .A(n2106), .B(n284), .Z(product[12]) );
  CIVXL U1783 ( .A(n1729), .Z(n1732) );
  CMXI2X1 U1784 ( .A0(n1731), .A1(n1086), .S(n1732), .Z(n815) );
  CIVX2 U1785 ( .A(n1087), .Z(n1734) );
  CIVX2 U1786 ( .A(n1730), .Z(n1735) );
  CENX1 U1787 ( .A(a[30]), .B(a[31]), .Z(n1730) );
  CENX1 U1788 ( .A(net183987), .B(a[30]), .Z(n1729) );
  CMXI2X1 U1789 ( .A0(n1088), .A1(n1733), .S(n1729), .Z(n799) );
  CND2XL U1790 ( .A(n1735), .B(n1734), .Z(n1731) );
  CENXL U1791 ( .A(net33076), .B(a[31]), .Z(n1087) );
  CENXL U1792 ( .A(net33422), .B(a[31]), .Z(n1086) );
  CENXL U1793 ( .A(n1783), .B(n1782), .Z(n1736) );
  CEO3XL U1794 ( .A(n735), .B(n733), .C(n726), .Z(n720) );
  CANR1XL U1795 ( .A(n269), .B(n278), .C(n1728), .Z(n1738) );
  COND2X1 U1796 ( .A(n1100), .B(n1812), .C(n1433), .D(n107), .Z(n801) );
  CND2X1 U1797 ( .A(n1764), .B(n1589), .Z(net178605) );
  CNR2X1 U1798 ( .A(n1764), .B(n1589), .Z(net179842) );
  CND2XL U1799 ( .A(n1753), .B(n1588), .Z(net33774) );
  CND2X1 U1800 ( .A(n1753), .B(n1758), .Z(net33776) );
  CENXL U1801 ( .A(n1793), .B(n1753), .Z(n1788) );
  CND2X1 U1802 ( .A(n566), .B(net171598), .Z(n1757) );
  CEOX1 U1803 ( .A(n665), .B(n650), .Z(n1739) );
  CND2X1 U1804 ( .A(n650), .B(n665), .Z(n1742) );
  CND3X1 U1805 ( .A(n1740), .B(n1741), .C(n1742), .Z(n643) );
  CNR2XL U1806 ( .A(n1148), .B(n82), .Z(n1743) );
  COR2X1 U1807 ( .A(n1743), .B(n1744), .Z(n805) );
  CIVXL U1808 ( .A(n2138), .Z(n1437) );
  CENX1 U1809 ( .A(n950), .B(n974), .Z(n1745) );
  CANR1X1 U1810 ( .A(n280), .B(n288), .C(n281), .Z(n279) );
  CEOXL U1811 ( .A(n1824), .B(n1669), .Z(n710) );
  CENXL U1812 ( .A(n1746), .B(n840), .Z(n508) );
  CENXL U1813 ( .A(n930), .B(n892), .Z(n1746) );
  CND2XL U1814 ( .A(n516), .B(n1761), .Z(net33755) );
  CND2XL U1815 ( .A(n1775), .B(n518), .Z(net33754) );
  CND2X1 U1816 ( .A(n1775), .B(net171496), .Z(net33752) );
  CIVX1 U1817 ( .A(n216), .Z(n342) );
  CND2XL U1818 ( .A(n231), .B(net178512), .Z(n224) );
  CIVXL U1819 ( .A(n167), .Z(n336) );
  CEOX1 U1820 ( .A(n440), .B(n463), .Z(n2119) );
  CFA1X1 U1821 ( .A(n968), .B(n1552), .CI(n992), .CO(n765), .S(n766) );
  CND2X2 U1822 ( .A(n1748), .B(n1749), .Z(n1750) );
  CND2X1 U1823 ( .A(n1874), .B(n1750), .Z(n1858) );
  CND2X2 U1824 ( .A(n1751), .B(n1752), .Z(product[11]) );
  CND2IX1 U1825 ( .B(a[24]), .A(n2169), .Z(n1975) );
  COND4CX4 U1826 ( .A(n1754), .B(n1755), .C(n1756), .D(n1757), .Z(n1753) );
  CIVX2 U1827 ( .A(net171595), .Z(n1765) );
  CIVX2 U1828 ( .A(net171604), .Z(n1766) );
  CIVX2 U1829 ( .A(net171598), .Z(n1755) );
  CIVX2 U1830 ( .A(net171596), .Z(n1768) );
  CNR2X2 U1831 ( .A(net171595), .B(net171594), .Z(n1770) );
  CIVX2 U1832 ( .A(net171602), .Z(n1771) );
  CNR2X2 U1833 ( .A(net171602), .B(net171600), .Z(n1772) );
  CIVX2 U1834 ( .A(net171593), .Z(n1773) );
  CIVX2 U1835 ( .A(net171472), .Z(n1774) );
  CENX2 U1836 ( .A(n1785), .B(n1765), .Z(n1756) );
  CMXI2X1 U1837 ( .A0(n1788), .A1(n1789), .S(n1588), .Z(n1764) );
  CEOX2 U1838 ( .A(n581), .B(n1583), .Z(net179820) );
  CND2IX1 U1839 ( .B(n1769), .A(n1795), .Z(n1777) );
  CIVX2 U1840 ( .A(net171592), .Z(n1783) );
  CND2IX1 U1841 ( .B(n1774), .A(n1786), .Z(n1796) );
  CIVX2 U1842 ( .A(n1753), .Z(n1797) );
  COND1X2 U1843 ( .A(n1767), .B(n1768), .C(n1798), .Z(n1795) );
  CIVX2 U1844 ( .A(n1795), .Z(n1784) );
  CND2X2 U1845 ( .A(net171595), .B(net171594), .Z(n1799) );
  COND1X2 U1846 ( .A(n1766), .B(n1770), .C(n1799), .Z(n1787) );
  COND1X2 U1847 ( .A(n1772), .B(n1773), .C(n1800), .Z(n1786) );
  CIVX2 U1848 ( .A(n1775), .Z(n1780) );
  CND2IX1 U1849 ( .B(n1774), .A(n1787), .Z(n1803) );
  CIVX2 U1850 ( .A(n1781), .Z(n1801) );
  CIVX2 U1851 ( .A(n1791), .Z(n560) );
  CENX2 U1852 ( .A(net171594), .B(net171604), .Z(n1785) );
  CEO3X2 U1853 ( .A(net171589), .B(n1784), .C(n1736), .Z(n1758) );
  CIVXL U1854 ( .A(net171589), .Z(n1769) );
  CENX2 U1855 ( .A(net171596), .B(net171597), .Z(n1804) );
  COND1X1 U1856 ( .A(n206), .B(n189), .C(n190), .Z(n188) );
  CANR1X2 U1857 ( .A(n187), .B(net179676), .C(n188), .Z(n186) );
  COR2X1 U1858 ( .A(net180312), .B(n512), .Z(n1805) );
  CANR1X1 U1859 ( .A(n1807), .B(net178507), .C(n212), .Z(n206) );
  CIVX2 U1860 ( .A(n214), .Z(n212) );
  CANR1XL U1861 ( .A(n1807), .B(net178507), .C(n212), .Z(net179529) );
  CND2X1 U1862 ( .A(n580), .B(n599), .Z(n217) );
  CND2X1 U1863 ( .A(net178605), .B(net180618), .Z(n189) );
  CNR2X1 U1864 ( .A(n205), .B(n189), .Z(n187) );
  CIVXL U1865 ( .A(net179842), .Z(net179838) );
  CND2X1 U1866 ( .A(n512), .B(net180312), .Z(n194) );
  CND2XL U1867 ( .A(net180618), .B(n194), .Z(n125) );
  CND3X1 U1868 ( .A(net33774), .B(net33775), .C(net33776), .Z(net180312) );
  COR2XL U1869 ( .A(net180312), .B(n512), .Z(net180618) );
  COR2X1 U1870 ( .A(n579), .B(n558), .Z(net178507) );
  CND2X1 U1871 ( .A(net178507), .B(n342), .Z(n205) );
  CND2XL U1872 ( .A(net178507), .B(n214), .Z(n127) );
  CND2X1 U1873 ( .A(n558), .B(n579), .Z(n214) );
  COND1XL U1874 ( .A(n158), .B(n186), .C(n159), .Z(n157) );
  CIVXL U1875 ( .A(n222), .Z(net179676) );
  CIVX2 U1876 ( .A(n223), .Z(n222) );
  CIVX2 U1877 ( .A(n229), .Z(n227) );
  COND2XL U1878 ( .A(n84), .B(n1144), .C(n82), .D(n1143), .Z(n866) );
  CFA1X1 U1879 ( .A(n862), .B(n826), .CI(n850), .CO(n509), .S(n510) );
  COND2X1 U1880 ( .A(n91), .B(n1127), .C(n89), .D(n1126), .Z(n850) );
  CIVXL U1881 ( .A(n712), .Z(n1809) );
  CIVX1 U1882 ( .A(n1809), .Z(n1810) );
  CNIVX2 U1883 ( .A(n846), .Z(n1811) );
  CENXL U1884 ( .A(a[26]), .B(n1835), .Z(net181698) );
  CENX1 U1885 ( .A(a[26]), .B(n1835), .Z(n1812) );
  CENXL U1886 ( .A(a[26]), .B(n2169), .Z(n105) );
  COAN1XL U1887 ( .A(n301), .B(n289), .C(n290), .Z(n1813) );
  CANR1X1 U1888 ( .A(n297), .B(n2018), .C(n292), .Z(n290) );
  COND1X1 U1889 ( .A(n325), .B(n323), .C(n324), .Z(n322) );
  CNR2IX1 U1890 ( .B(net33078), .A(n24), .Z(n1024) );
  CND2IX2 U1891 ( .B(n1591), .A(n185), .Z(n1998) );
  CNR2X2 U1892 ( .A(n1664), .B(n511), .Z(n183) );
  CENX2 U1893 ( .A(a[10]), .B(n2202), .Z(n1416) );
  COND2XL U1894 ( .A(n97), .B(n1113), .C(n95), .D(n1112), .Z(n837) );
  CIVXL U1895 ( .A(n58), .Z(net180673) );
  CIVX1 U1896 ( .A(net180673), .Z(net180674) );
  CEOX2 U1897 ( .A(n458), .B(n454), .Z(n1944) );
  COAN1X1 U1898 ( .A(n255), .B(n251), .C(n252), .Z(n248) );
  CND2X1 U1899 ( .A(n2034), .B(n2032), .Z(n255) );
  CND2X1 U1900 ( .A(n672), .B(n2035), .Z(n252) );
  CENX1 U1901 ( .A(n2193), .B(a[10]), .Z(n1815) );
  CENX1 U1902 ( .A(n2193), .B(a[10]), .Z(n1816) );
  CND2X1 U1903 ( .A(n629), .B(n612), .Z(n1817) );
  CND2XL U1904 ( .A(n629), .B(n614), .Z(n1818) );
  CND2X1 U1905 ( .A(n612), .B(n614), .Z(n1819) );
  CND3X2 U1906 ( .A(n1817), .B(n1818), .C(n1819), .Z(n605) );
  CEOX2 U1907 ( .A(n590), .B(n607), .Z(n1820) );
  CEOX2 U1908 ( .A(n1820), .B(n605), .Z(n584) );
  CND2XL U1909 ( .A(n607), .B(n590), .Z(n1821) );
  CND2XL U1910 ( .A(n590), .B(n605), .Z(n1822) );
  CND2XL U1911 ( .A(n607), .B(n605), .Z(n1823) );
  CND3XL U1912 ( .A(n1821), .B(n1822), .C(n1823), .Z(n583) );
  CHA1X1 U1913 ( .A(n847), .B(n873), .CO(n433), .S(n434) );
  COND2X1 U1914 ( .A(n91), .B(n1124), .C(n89), .D(n1123), .Z(n847) );
  CEOX1 U1915 ( .A(n1041), .B(n987), .Z(n1824) );
  CND2XL U1916 ( .A(n987), .B(n1041), .Z(n1827) );
  COND2XL U1917 ( .A(n18), .B(n1327), .C(n1326), .D(n15), .Z(n1041) );
  CENX1 U1918 ( .A(net33422), .B(n2203), .Z(n1203) );
  CND2X2 U1919 ( .A(n1415), .B(n58), .Z(n61) );
  CEO3X2 U1920 ( .A(n996), .B(n1022), .C(n1050), .Z(n790) );
  CEOX1 U1921 ( .A(n1080), .B(n793), .Z(n1828) );
  CEOX2 U1922 ( .A(n1828), .B(n790), .Z(n788) );
  CND2XL U1923 ( .A(n996), .B(n1022), .Z(n1829) );
  CND2X1 U1924 ( .A(n996), .B(n1050), .Z(n1830) );
  CND2XL U1925 ( .A(n1022), .B(n1050), .Z(n1831) );
  CND3X1 U1926 ( .A(n1829), .B(n1830), .C(n1831), .Z(n789) );
  CND2X1 U1927 ( .A(n1080), .B(n793), .Z(n1832) );
  CND2XL U1928 ( .A(n1080), .B(n790), .Z(n1833) );
  CND2XL U1929 ( .A(n793), .B(n790), .Z(n1834) );
  CND3X1 U1930 ( .A(n1832), .B(n1833), .C(n1834), .Z(n787) );
  CNIVX4 U1931 ( .A(n99), .Z(n1835) );
  CND2XL U1932 ( .A(n828), .B(n872), .Z(n1886) );
  CND2XL U1933 ( .A(n828), .B(n926), .Z(n1887) );
  COND2X1 U1934 ( .A(n91), .B(n1131), .C(n89), .D(n1130), .Z(n854) );
  COND2XL U1935 ( .A(n91), .B(n1123), .C(n89), .D(n1122), .Z(n846) );
  CND2X4 U1936 ( .A(n1416), .B(n50), .Z(n2117) );
  CNIVX4 U1937 ( .A(n93), .Z(n1933) );
  CND2X1 U1938 ( .A(n1662), .B(n131), .Z(n1996) );
  CIVX2 U1939 ( .A(n2169), .Z(n1973) );
  COND2X1 U1940 ( .A(n61), .B(n1691), .C(n58), .D(n1205), .Z(n808) );
  COND2X1 U1941 ( .A(n1114), .B(n97), .C(n95), .D(n1113), .Z(n838) );
  CND2IXL U1942 ( .B(n129), .A(n230), .Z(n1994) );
  CEOX1 U1943 ( .A(n957), .B(n881), .Z(n1836) );
  CEOX2 U1944 ( .A(n1836), .B(n1607), .Z(n616) );
  CND2XL U1945 ( .A(n804), .B(n881), .Z(n1837) );
  CND2XL U1946 ( .A(n957), .B(n804), .Z(n1838) );
  CND2XL U1947 ( .A(n881), .B(n957), .Z(n1839) );
  CND3X1 U1948 ( .A(n1837), .B(n1838), .C(n1839), .Z(n615) );
  COND2XL U1949 ( .A(n44), .B(n1240), .C(n1239), .D(n42), .Z(n957) );
  CND2XL U1950 ( .A(n615), .B(n613), .Z(n1890) );
  CND2X1 U1951 ( .A(n721), .B(n723), .Z(n1882) );
  CND2X1 U1952 ( .A(n712), .B(n721), .Z(n1880) );
  CND2X1 U1953 ( .A(n831), .B(n975), .Z(n1840) );
  CND2X1 U1954 ( .A(n831), .B(n951), .Z(n1841) );
  CND2X1 U1955 ( .A(n975), .B(n951), .Z(n1842) );
  CND3X1 U1956 ( .A(n1840), .B(n1841), .C(n1842), .Z(n479) );
  COR2X1 U1957 ( .A(n1106), .B(n1747), .Z(n1843) );
  CND2X2 U1958 ( .A(n1843), .B(n1844), .Z(n831) );
  COND2XL U1959 ( .A(n44), .B(n1234), .C(n1233), .D(n42), .Z(n951) );
  CND2X1 U1960 ( .A(n1934), .B(n1672), .Z(n1937) );
  CENXL U1961 ( .A(n2171), .B(b[24]), .Z(n1315) );
  CENXL U1962 ( .A(n2171), .B(n1384), .Z(n1318) );
  CENXL U1963 ( .A(n2171), .B(n1387), .Z(n1321) );
  CENXL U1964 ( .A(n2171), .B(n2157), .Z(n1331) );
  CND2IXL U1965 ( .B(net33078), .A(n2171), .Z(n1340) );
  CIVX1 U1966 ( .A(net184424), .Z(net179546) );
  CENX1 U1967 ( .A(n479), .B(n477), .Z(n1845) );
  CND2X1 U1968 ( .A(n719), .B(n1846), .Z(n1849) );
  CND2X2 U1969 ( .A(n1848), .B(n1849), .Z(n1900) );
  CIVXL U1970 ( .A(n710), .Z(n1846) );
  CND2X2 U1971 ( .A(n1984), .B(n1985), .Z(n855) );
  CND2X1 U1972 ( .A(n1411), .B(n1962), .Z(n1984) );
  CND2XL U1973 ( .A(n429), .B(n425), .Z(n1850) );
  CND2XL U1974 ( .A(n429), .B(n427), .Z(n1851) );
  CND2XL U1975 ( .A(n425), .B(n427), .Z(n1852) );
  CND3XL U1976 ( .A(n1850), .B(n1851), .C(n1852), .Z(n393) );
  COND2X1 U1977 ( .A(n36), .B(n1276), .C(n1275), .D(net178746), .Z(n992) );
  CND2XL U1978 ( .A(n898), .B(n916), .Z(n2141) );
  CND2XL U1979 ( .A(n832), .B(n1602), .Z(n1853) );
  CND2XL U1980 ( .A(n832), .B(n952), .Z(n1854) );
  CND2XL U1981 ( .A(n1602), .B(n952), .Z(n1855) );
  CND3X1 U1982 ( .A(n1853), .B(n1854), .C(n1855), .Z(n505) );
  COND2XL U1983 ( .A(n44), .B(n1235), .C(n1234), .D(n42), .Z(n952) );
  CND2XL U1984 ( .A(n567), .B(n569), .Z(n2148) );
  CND2XL U1985 ( .A(n548), .B(n567), .Z(n2146) );
  CNIVX3 U1986 ( .A(n63), .Z(n1857) );
  CNR2IX1 U1987 ( .B(n89), .A(n1132), .Z(n1962) );
  CEOX2 U1988 ( .A(a[18]), .B(n2167), .Z(n1412) );
  CEOX2 U1989 ( .A(n2038), .B(n2039), .Z(n1859) );
  CEOX2 U1990 ( .A(n1859), .B(n2040), .Z(n656) );
  CND2XL U1991 ( .A(n2040), .B(n2039), .Z(n1860) );
  CND2XL U1992 ( .A(n2040), .B(n2038), .Z(n1861) );
  CND2XL U1993 ( .A(n2039), .B(n2038), .Z(n1862) );
  CND3XL U1994 ( .A(n1860), .B(n1861), .C(n1862), .Z(n655) );
  CIVXL U1995 ( .A(n1439), .Z(n1863) );
  COND2X1 U1996 ( .A(n27), .B(n1306), .C(n1305), .D(n24), .Z(n1021) );
  COND2X1 U1997 ( .A(n27), .B(n1303), .C(n1302), .D(n24), .Z(n1018) );
  COND2X1 U1998 ( .A(n27), .B(n1302), .C(n1301), .D(n24), .Z(n1017) );
  CND2IX4 U1999 ( .B(n2011), .A(n24), .Z(n27) );
  CHA1X1 U2000 ( .A(n945), .B(n809), .CO(n757), .S(n758) );
  COND2X1 U2001 ( .A(n2117), .B(n1654), .C(n1816), .D(n1228), .Z(n809) );
  CEOX1 U2002 ( .A(n631), .B(n633), .Z(n1864) );
  CND2X1 U2003 ( .A(n616), .B(n633), .Z(n1865) );
  CND2X1 U2004 ( .A(n616), .B(n631), .Z(n1866) );
  CND2X1 U2005 ( .A(n633), .B(n631), .Z(n1867) );
  CND3X1 U2006 ( .A(n1865), .B(n1866), .C(n1867), .Z(n607) );
  CFA1XL U2007 ( .A(n936), .B(n1066), .CI(n1008), .CO(n631), .S(n632) );
  CND3X1 U2008 ( .A(net180364), .B(net180365), .C(net180366), .Z(n429) );
  CENXL U2009 ( .A(n2152), .B(n1623), .Z(n1096) );
  CND2XL U2010 ( .A(n840), .B(n892), .Z(n1868) );
  CND2XL U2011 ( .A(n840), .B(n930), .Z(n1869) );
  CND2X1 U2012 ( .A(n892), .B(n930), .Z(n1870) );
  CND3X1 U2013 ( .A(n1868), .B(n1869), .C(n1870), .Z(n507) );
  CENX4 U2014 ( .A(n2166), .B(a[18]), .Z(n82) );
  CND2XL U2015 ( .A(n948), .B(n822), .Z(n1871) );
  CND2X1 U2016 ( .A(n948), .B(n888), .Z(n1872) );
  CND2XL U2017 ( .A(n822), .B(n888), .Z(n1873) );
  CND3X1 U2018 ( .A(n1871), .B(n1872), .C(n1873), .Z(n399) );
  CND2XL U2019 ( .A(n406), .B(n404), .Z(n1874) );
  CND2XL U2020 ( .A(n1576), .B(n400), .Z(n1875) );
  CND2XL U2021 ( .A(n404), .B(n400), .Z(n1876) );
  CND3XL U2022 ( .A(n1615), .B(n1875), .C(n1876), .Z(n391) );
  CIVX2 U2023 ( .A(n39), .Z(n2199) );
  CFA1X1 U2024 ( .A(n856), .B(n1550), .CI(n868), .CO(n635), .S(n636) );
  CNR2IX1 U2025 ( .B(net33078), .A(n89), .Z(n856) );
  CEOX2 U2026 ( .A(n723), .B(n721), .Z(n1879) );
  CEOX2 U2027 ( .A(n1879), .B(n1810), .Z(n706) );
  CND2X1 U2028 ( .A(n712), .B(n723), .Z(n1881) );
  CND3X1 U2029 ( .A(n1880), .B(n1881), .C(n1882), .Z(n705) );
  COR2X1 U2030 ( .A(n1695), .B(n61), .Z(n1883) );
  CND2X2 U2031 ( .A(n1883), .B(n1884), .Z(n921) );
  CFA1XL U2032 ( .A(n964), .B(n1072), .CI(n1042), .CO(n723), .S(n724) );
  CEOX1 U2033 ( .A(n926), .B(n872), .Z(n1885) );
  CEOX1 U2034 ( .A(n1885), .B(n828), .Z(n404) );
  CND2X1 U2035 ( .A(n872), .B(n926), .Z(n1888) );
  CND3XL U2036 ( .A(n1886), .B(n1887), .C(n1888), .Z(n403) );
  CEO3X1 U2037 ( .A(n405), .B(n403), .C(n399), .Z(n372) );
  CFA1X1 U2038 ( .A(n955), .B(n853), .CI(n879), .CO(n575), .S(n576) );
  COND2X1 U2039 ( .A(n91), .B(n1130), .C(n89), .D(n1129), .Z(n853) );
  CND2XL U2040 ( .A(n829), .B(n889), .Z(n1907) );
  CND2XL U2041 ( .A(n829), .B(n949), .Z(n1908) );
  CND2XL U2042 ( .A(n841), .B(n802), .Z(n1896) );
  CND2X2 U2043 ( .A(n2014), .B(n2015), .Z(product[31]) );
  CND2XL U2044 ( .A(n615), .B(n617), .Z(n1889) );
  CND2XL U2045 ( .A(n617), .B(n613), .Z(n1891) );
  CND3XL U2046 ( .A(n1889), .B(n1890), .C(n1891), .Z(n589) );
  CND2XL U2047 ( .A(n460), .B(n477), .Z(n1892) );
  CND2XL U2048 ( .A(n460), .B(n479), .Z(n1893) );
  CND2XL U2049 ( .A(n477), .B(n479), .Z(n1894) );
  CND3XL U2050 ( .A(n1892), .B(n1893), .C(n1894), .Z(n447) );
  CIVXL U2051 ( .A(net179838), .Z(net180217) );
  COR2X1 U2052 ( .A(n89), .B(n1131), .Z(n1985) );
  CND2IX2 U2053 ( .B(n2006), .A(n95), .Z(n97) );
  CENXL U2054 ( .A(n532), .B(n1895), .Z(n2132) );
  CFA1X1 U2055 ( .A(n864), .B(n1666), .CI(n834), .CO(n555), .S(n556) );
  CND2X2 U2056 ( .A(n488), .B(n511), .Z(n184) );
  CND2XL U2057 ( .A(n824), .B(n950), .Z(n1911) );
  CND2XL U2058 ( .A(n824), .B(n974), .Z(n1910) );
  CIVXL U2059 ( .A(n1835), .Z(n1434) );
  CND2X2 U2060 ( .A(n351), .B(n2107), .Z(n137) );
  CIVX3 U2061 ( .A(n2108), .Z(n351) );
  CENX1 U2062 ( .A(n2151), .B(n2203), .Z(n1202) );
  CNR2X1 U2063 ( .A(n716), .B(n727), .Z(n271) );
  COND2X1 U2064 ( .A(net179858), .B(n1090), .C(n1089), .D(n110), .Z(n817) );
  CND2X1 U2065 ( .A(n841), .B(n953), .Z(n1897) );
  CNIVX2 U2066 ( .A(n841), .Z(n1899) );
  COND2XL U2067 ( .A(n44), .B(n1236), .C(n1235), .D(n42), .Z(n953) );
  CEO3X2 U2068 ( .A(n1013), .B(n714), .C(n725), .Z(n708) );
  CND2X1 U2069 ( .A(n1013), .B(n714), .Z(n1901) );
  CND2X1 U2070 ( .A(n1013), .B(n725), .Z(n1902) );
  CND2X1 U2071 ( .A(n714), .B(n725), .Z(n1903) );
  CND3X2 U2072 ( .A(n1901), .B(n1902), .C(n1903), .Z(n707) );
  CND2XL U2073 ( .A(n719), .B(n710), .Z(n1904) );
  CND2XL U2074 ( .A(n719), .B(n708), .Z(n1906) );
  CND3X1 U2075 ( .A(n1904), .B(n1905), .C(n1906), .Z(n703) );
  CEOX1 U2076 ( .A(n949), .B(n889), .Z(net180068) );
  CND2X1 U2077 ( .A(n889), .B(n949), .Z(n1909) );
  CND2X1 U2078 ( .A(n974), .B(n950), .Z(n1912) );
  COND2XL U2079 ( .A(n44), .B(n1233), .C(n1232), .D(n42), .Z(n950) );
  CEOX1 U2080 ( .A(n2045), .B(n2047), .Z(n1913) );
  CEOX2 U2081 ( .A(n1913), .B(n622), .Z(n620) );
  CND2XL U2082 ( .A(n622), .B(n2047), .Z(n1914) );
  CND2XL U2083 ( .A(n622), .B(n2045), .Z(n1915) );
  CND2XL U2084 ( .A(n2047), .B(n2045), .Z(n1916) );
  CND3XL U2085 ( .A(n1914), .B(n1915), .C(n1916), .Z(n619) );
  CND2XL U2086 ( .A(n246), .B(n132), .Z(n1919) );
  CND2X1 U2087 ( .A(n1917), .B(n1918), .Z(n1920) );
  CIVXL U2088 ( .A(n246), .Z(n1917) );
  CIVXL U2089 ( .A(n132), .Z(n1918) );
  CND2X1 U2090 ( .A(n346), .B(n245), .Z(n132) );
  CENXL U2091 ( .A(n2008), .B(n548), .Z(n542) );
  CIVX1 U2092 ( .A(a[22]), .Z(n1981) );
  CENX1 U2093 ( .A(n2205), .B(a[12]), .Z(n1415) );
  CHA1X1 U2094 ( .A(n808), .B(n965), .CO(n737), .S(n738) );
  CND2X1 U2095 ( .A(n2002), .B(n2003), .Z(product[15]) );
  CND2XL U2096 ( .A(n858), .B(n818), .Z(n1921) );
  CND2X1 U2097 ( .A(n858), .B(n906), .Z(n1922) );
  CND2XL U2098 ( .A(n818), .B(n906), .Z(n1923) );
  CND2XL U2099 ( .A(n423), .B(n398), .Z(n1924) );
  CND2XL U2100 ( .A(n423), .B(n402), .Z(n1925) );
  CND2XL U2101 ( .A(n398), .B(n402), .Z(n1926) );
  CND3XL U2102 ( .A(n1924), .B(n1925), .C(n1926), .Z(n389) );
  COR2XL U2103 ( .A(n1090), .B(net184424), .Z(n1927) );
  CENX2 U2104 ( .A(n123), .B(n2000), .Z(product[27]) );
  CND2X2 U2105 ( .A(n1998), .B(n1999), .Z(n2000) );
  CNIVX4 U2106 ( .A(n86), .Z(n1928) );
  CENXL U2107 ( .A(n2163), .B(n2204), .Z(n1190) );
  CENXL U2108 ( .A(n2160), .B(n2204), .Z(n1193) );
  CENXL U2109 ( .A(n2161), .B(n2204), .Z(n1192) );
  CENXL U2110 ( .A(n2162), .B(n2204), .Z(n1191) );
  CENXL U2111 ( .A(n2159), .B(n2204), .Z(n1194) );
  CENXL U2112 ( .A(n2156), .B(n2204), .Z(n1197) );
  CENXL U2113 ( .A(n2158), .B(n2204), .Z(n1195) );
  CENXL U2114 ( .A(n2157), .B(n2204), .Z(n1196) );
  CND2XL U2115 ( .A(n733), .B(n726), .Z(n1929) );
  CND2XL U2116 ( .A(n733), .B(n735), .Z(n1930) );
  CND2XL U2117 ( .A(n726), .B(n735), .Z(n1931) );
  CND3X1 U2118 ( .A(n1929), .B(n1930), .C(n1931), .Z(n719) );
  CFA1XL U2119 ( .A(n943), .B(n1073), .CI(n1015), .CO(n735), .S(n736) );
  CFA1XL U2120 ( .A(n989), .B(n923), .CI(n1043), .CO(n733), .S(n734) );
  CND2IX2 U2121 ( .B(n2026), .A(n66), .Z(n1932) );
  CND2XL U2122 ( .A(a[16]), .B(n1935), .Z(n1936) );
  CIVXL U2123 ( .A(a[16]), .Z(n1934) );
  CNIVX4 U2124 ( .A(n71), .Z(n2166) );
  CIVXL U2125 ( .A(n1933), .Z(n1435) );
  CND2X1 U2126 ( .A(n347), .B(n252), .Z(n133) );
  CENX1 U2127 ( .A(n1963), .B(n171), .Z(product[28]) );
  CEO3XL U2128 ( .A(n2118), .B(n1547), .C(n800), .Z(n432) );
  CND2XL U2129 ( .A(n453), .B(n451), .Z(n1941) );
  CND2XL U2130 ( .A(n432), .B(n453), .Z(n1942) );
  CND2XL U2131 ( .A(n432), .B(n451), .Z(n1943) );
  CND3XL U2132 ( .A(n1943), .B(n1942), .C(n1941), .Z(n419) );
  CND2XL U2133 ( .A(n456), .B(n454), .Z(n1945) );
  CND2XL U2134 ( .A(n456), .B(n458), .Z(n1946) );
  CND2XL U2135 ( .A(n454), .B(n458), .Z(n1947) );
  CND3XL U2136 ( .A(n1945), .B(n1946), .C(n1947), .Z(n445) );
  CFA1XL U2137 ( .A(n860), .B(n928), .CI(n874), .CO(n457), .S(n458) );
  CNR2X2 U2138 ( .A(n408), .B(n435), .Z(n1986) );
  CND2X1 U2139 ( .A(n467), .B(n469), .Z(n1956) );
  CND2X1 U2140 ( .A(n2080), .B(n467), .Z(n1954) );
  CENX2 U2141 ( .A(a[14]), .B(n2165), .Z(n2026) );
  CENXL U2142 ( .A(net33076), .B(n1835), .Z(n1108) );
  CENXL U2143 ( .A(n2156), .B(n1835), .Z(n1101) );
  CND2IXL U2144 ( .B(net33078), .A(n1835), .Z(n1109) );
  CENXL U2145 ( .A(n2151), .B(n1835), .Z(n1106) );
  CENXL U2146 ( .A(n2155), .B(n1835), .Z(n1102) );
  CENXL U2147 ( .A(n2154), .B(n1835), .Z(n1103) );
  CENXL U2148 ( .A(n2153), .B(n2169), .Z(n1104) );
  CNR2X2 U2149 ( .A(n1610), .B(n183), .Z(n172) );
  COND2X1 U2150 ( .A(n1117), .B(n97), .C(n95), .D(n1116), .Z(n841) );
  CND2X1 U2151 ( .A(net171496), .B(n518), .Z(n2149) );
  CEOX2 U2152 ( .A(net179820), .B(n560), .Z(n558) );
  CEO3X2 U2153 ( .A(n2067), .B(n2062), .C(n2068), .Z(n470) );
  CND2XL U2154 ( .A(n2067), .B(n2062), .Z(n1950) );
  CND2XL U2155 ( .A(n2067), .B(n2068), .Z(n1951) );
  CND2X1 U2156 ( .A(n2062), .B(n2068), .Z(n1952) );
  CND3X1 U2157 ( .A(n1950), .B(n1951), .C(n1952), .Z(n469) );
  CND2X1 U2158 ( .A(n2080), .B(n469), .Z(n1955) );
  CND3X2 U2159 ( .A(n1954), .B(n1955), .C(n1956), .Z(n439) );
  CANR1XL U2160 ( .A(n1682), .B(n1558), .C(n161), .Z(n1957) );
  CND3X1 U2161 ( .A(n2123), .B(n2124), .C(n2125), .Z(n435) );
  CNR2X1 U2162 ( .A(n1986), .B(n167), .Z(n160) );
  COND2X1 U2163 ( .A(n1120), .B(n95), .C(n1435), .D(n97), .Z(n803) );
  CND2X1 U2164 ( .A(n1677), .B(n120), .Z(n1988) );
  COND2XL U2165 ( .A(n36), .B(n1262), .C(n1261), .D(net178746), .Z(n978) );
  COND2XL U2166 ( .A(n36), .B(n1260), .C(n1259), .D(net178746), .Z(n976) );
  COND2XL U2167 ( .A(n36), .B(n1261), .C(n1260), .D(net178746), .Z(n977) );
  COND2XL U2168 ( .A(n36), .B(n1264), .C(n1263), .D(net178746), .Z(n980) );
  COND2XL U2169 ( .A(n36), .B(n1265), .C(n1264), .D(net178746), .Z(n981) );
  COND2XL U2170 ( .A(n36), .B(n1270), .C(n1269), .D(net178746), .Z(n986) );
  COND2XL U2171 ( .A(n36), .B(n1271), .C(n1270), .D(net178746), .Z(n987) );
  COND2XL U2172 ( .A(n2117), .B(n1212), .C(n1211), .D(n1816), .Z(n930) );
  COND2XL U2173 ( .A(n2117), .B(n1217), .C(n1216), .D(n1816), .Z(n935) );
  COND2X1 U2174 ( .A(n1227), .B(n2117), .C(n1815), .D(n1226), .Z(n945) );
  CANR1XL U2175 ( .A(n314), .B(n2022), .C(n311), .Z(n1959) );
  CIVX2 U2176 ( .A(n313), .Z(n311) );
  CFA1X1 U2177 ( .A(n924), .B(n966), .CI(n944), .CO(n747), .S(n748) );
  CEN3X1 U2178 ( .A(n1960), .B(n374), .C(n395), .Z(n369) );
  CEN3X2 U2179 ( .A(n971), .B(n997), .C(n1025), .Z(n1960) );
  CNIVX4 U2180 ( .A(n79), .Z(n2138) );
  CENXL U2181 ( .A(n2164), .B(n1672), .Z(n1149) );
  CENXL U2182 ( .A(n2157), .B(n1672), .Z(n1156) );
  CENXL U2183 ( .A(n2159), .B(n1672), .Z(n1154) );
  CENXL U2184 ( .A(n2163), .B(n1672), .Z(n1150) );
  CENXL U2185 ( .A(n2162), .B(n1672), .Z(n1151) );
  CENXL U2186 ( .A(n2158), .B(n1672), .Z(n1155) );
  CENXL U2187 ( .A(n2161), .B(n1672), .Z(n1152) );
  CENXL U2188 ( .A(n2160), .B(n1672), .Z(n1153) );
  CENXL U2189 ( .A(n2156), .B(n1672), .Z(n1157) );
  CENXL U2190 ( .A(net33078), .B(n1672), .Z(n1164) );
  CENXL U2191 ( .A(n2155), .B(n1672), .Z(n1158) );
  CENXL U2192 ( .A(n2154), .B(n1672), .Z(n1159) );
  CENXL U2193 ( .A(net33422), .B(n1672), .Z(n1163) );
  CENXL U2194 ( .A(n2152), .B(n1672), .Z(n1161) );
  CENXL U2195 ( .A(n2153), .B(n1672), .Z(n1160) );
  CENXL U2196 ( .A(n2151), .B(n1672), .Z(n1162) );
  CANR1X1 U2197 ( .A(n231), .B(n1661), .C(n232), .Z(n230) );
  CIVX4 U2198 ( .A(n2205), .Z(n2203) );
  CFA1X1 U2199 ( .A(n2036), .B(n2037), .CI(n2033), .S(n1961) );
  CNR2X1 U2200 ( .A(n2110), .B(n2108), .Z(n269) );
  CENXL U2201 ( .A(n2162), .B(n2138), .Z(n1134) );
  CENXL U2202 ( .A(n2154), .B(n2138), .Z(n1142) );
  CENXL U2203 ( .A(n2153), .B(n2138), .Z(n1143) );
  CENXL U2204 ( .A(n2157), .B(n2138), .Z(n1139) );
  CENXL U2205 ( .A(net33076), .B(n2138), .Z(n1147) );
  CENXL U2206 ( .A(n2155), .B(n2138), .Z(n1141) );
  CENXL U2207 ( .A(n2156), .B(n2138), .Z(n1140) );
  CENXL U2208 ( .A(n2159), .B(n2138), .Z(n1137) );
  CENXL U2209 ( .A(n2158), .B(n2138), .Z(n1138) );
  CENXL U2210 ( .A(n2152), .B(n2138), .Z(n1144) );
  CENXL U2211 ( .A(n2151), .B(n2138), .Z(n1145) );
  CND2IXL U2212 ( .B(net33078), .A(n2138), .Z(n1148) );
  COND2X1 U2213 ( .A(n1697), .B(n1164), .C(n74), .D(n1163), .Z(n885) );
  CANR1X1 U2214 ( .A(n2019), .B(n300), .C(n297), .Z(n295) );
  CND2X4 U2215 ( .A(n1982), .B(n1983), .Z(n95) );
  CND2X1 U2216 ( .A(a[22]), .B(n2168), .Z(n1982) );
  COND1X1 U2217 ( .A(n2105), .B(n2113), .C(n2104), .Z(n284) );
  CENXL U2218 ( .A(n142), .B(n306), .Z(product[8]) );
  CEO3X1 U2219 ( .A(n925), .B(n817), .C(n827), .Z(n376) );
  CIVX4 U2220 ( .A(n48), .Z(n2202) );
  CFA1X1 U2221 ( .A(n954), .B(n842), .CI(n894), .CO(n553), .S(n554) );
  CFA1X1 U2222 ( .A(n534), .B(n553), .CI(n555), .CO(n523), .S(n524) );
  CND2X2 U2223 ( .A(n1408), .B(n1812), .Z(n107) );
  CENXL U2224 ( .A(n2200), .B(n1384), .Z(n1206) );
  COND2XL U2225 ( .A(n61), .B(n1192), .C(n1191), .D(net180674), .Z(n911) );
  CENXL U2226 ( .A(n2200), .B(n2162), .Z(n1214) );
  CENXL U2227 ( .A(n2200), .B(n1389), .Z(n1211) );
  CENXL U2228 ( .A(n2200), .B(n2163), .Z(n1213) );
  CENXL U2229 ( .A(n2200), .B(n1387), .Z(n1209) );
  CENXL U2230 ( .A(n2200), .B(n1388), .Z(n1210) );
  CENXL U2231 ( .A(n2200), .B(n1386), .Z(n1208) );
  CENXL U2232 ( .A(n2200), .B(n2164), .Z(n1212) );
  CENXL U2233 ( .A(n2200), .B(n1385), .Z(n1207) );
  COND2XL U2234 ( .A(n61), .B(n1196), .C(n58), .D(n1195), .Z(n915) );
  CENXL U2235 ( .A(n2200), .B(n2161), .Z(n1215) );
  COND2XL U2236 ( .A(n61), .B(n1199), .C(n58), .D(n1198), .Z(n918) );
  CENXL U2237 ( .A(n2200), .B(n2160), .Z(n1216) );
  COND2XL U2238 ( .A(n1204), .B(n61), .C(n58), .D(n1203), .Z(n923) );
  CENXL U2239 ( .A(n2200), .B(n2159), .Z(n1217) );
  CENXL U2240 ( .A(n2156), .B(n2200), .Z(n1220) );
  CNR2IX1 U2241 ( .B(net33078), .A(n58), .Z(n924) );
  CAN2XL U2242 ( .A(n336), .B(n170), .Z(n1963) );
  CENXL U2243 ( .A(n2154), .B(net182741), .Z(n1094) );
  CENXL U2244 ( .A(net180562), .B(net33076), .Z(n1099) );
  CND2IXL U2245 ( .B(net33078), .A(net182741), .Z(n1100) );
  CENX2 U2246 ( .A(a[16]), .B(n1856), .Z(n74) );
  CND2IXL U2247 ( .B(net33078), .A(net183987), .Z(n1093) );
  CIVXL U2248 ( .A(net183987), .Z(n1432) );
  CENXL U2249 ( .A(n1696), .B(n1386), .Z(n1185) );
  CENXL U2250 ( .A(n2164), .B(n1696), .Z(n1189) );
  CENXL U2251 ( .A(n1696), .B(n1389), .Z(n1188) );
  CENXL U2252 ( .A(n2153), .B(n2203), .Z(n1200) );
  CENXL U2253 ( .A(n2155), .B(n2203), .Z(n1198) );
  CENXL U2254 ( .A(n2154), .B(n2203), .Z(n1199) );
  CND2IX1 U2255 ( .B(n157), .A(n1987), .Z(n1989) );
  COND1X1 U2256 ( .A(n2110), .B(n2107), .C(n2109), .Z(n1964) );
  CND2IX1 U2257 ( .B(n268), .A(n2010), .Z(n2003) );
  COND1XL U2258 ( .A(n2107), .B(n2110), .C(n2109), .Z(n270) );
  CANR1X1 U2259 ( .A(n269), .B(n278), .C(n1964), .Z(n268) );
  CENXL U2260 ( .A(n2157), .B(n2200), .Z(n1219) );
  CENXL U2261 ( .A(n2158), .B(n2200), .Z(n1218) );
  CENXL U2262 ( .A(n2155), .B(n2201), .Z(n1221) );
  CENXL U2263 ( .A(n2154), .B(n2201), .Z(n1222) );
  CENXL U2264 ( .A(n2153), .B(n2201), .Z(n1223) );
  CND2IXL U2265 ( .B(net33078), .A(n2201), .Z(n1228) );
  CENXL U2266 ( .A(n2152), .B(n2201), .Z(n1224) );
  CENXL U2267 ( .A(net33076), .B(n2201), .Z(n1227) );
  CNIVX2 U2268 ( .A(n900), .Z(n1965) );
  COND2XL U2269 ( .A(n84), .B(n1138), .C(n82), .D(n1137), .Z(n860) );
  COND2XL U2270 ( .A(n84), .B(n1136), .C(n82), .D(n1135), .Z(n858) );
  COND2XL U2271 ( .A(n84), .B(n1139), .C(n82), .D(n1138), .Z(n861) );
  COND2XL U2272 ( .A(n84), .B(n1141), .C(n82), .D(n1140), .Z(n863) );
  COND2XL U2273 ( .A(n1102), .B(n1747), .C(n1814), .D(n1101), .Z(n827) );
  CENXL U2274 ( .A(n125), .B(n195), .Z(product[25]) );
  CIVX2 U2275 ( .A(n173), .Z(n175) );
  CENXL U2276 ( .A(net33078), .B(n2204), .Z(n1204) );
  CND2IX2 U2277 ( .B(n2016), .A(n1726), .Z(n1991) );
  CIVX1 U2278 ( .A(n899), .Z(n1966) );
  CIVX2 U2279 ( .A(n1966), .Z(n1967) );
  CFA1X1 U2280 ( .A(n573), .B(n556), .CI(n571), .CO(n545), .S(n546) );
  CIVX1 U2281 ( .A(n120), .Z(n1987) );
  CENXL U2282 ( .A(n124), .B(n185), .Z(product[26]) );
  CANR1X1 U2283 ( .A(n172), .B(net179617), .C(n1609), .Z(n171) );
  CNR2X1 U2284 ( .A(n702), .B(n715), .Z(n266) );
  COND2XL U2285 ( .A(n1570), .B(n1180), .C(n66), .D(n1179), .Z(n900) );
  COND2XL U2286 ( .A(n1570), .B(n1179), .C(n66), .D(n1178), .Z(n899) );
  CNR2IX1 U2287 ( .B(net33078), .A(n82), .Z(n870) );
  CIVX1 U2288 ( .A(n2111), .Z(n265) );
  CEOX2 U2289 ( .A(net180562), .B(a[26]), .Z(n1408) );
  CEO3XL U2290 ( .A(n947), .B(n1055), .C(n815), .Z(n374) );
  CIVX2 U2291 ( .A(n244), .Z(n346) );
  CNR2X2 U2292 ( .A(n656), .B(n671), .Z(n244) );
  CND2IXL U2293 ( .B(net33078), .A(n1933), .Z(n1120) );
  CENXL U2294 ( .A(net33076), .B(n1933), .Z(n1119) );
  CENXL U2295 ( .A(net33422), .B(n1933), .Z(n1118) );
  CENXL U2296 ( .A(n2158), .B(n1933), .Z(n1110) );
  CENXL U2297 ( .A(n2152), .B(n1933), .Z(n1116) );
  CENXL U2298 ( .A(n2153), .B(n1933), .Z(n1115) );
  CENXL U2299 ( .A(n2151), .B(n1933), .Z(n1117) );
  CENXL U2300 ( .A(n2154), .B(n1933), .Z(n1114) );
  COND2XL U2301 ( .A(n91), .B(n1125), .C(n89), .D(n1124), .Z(n848) );
  CEO3X1 U2302 ( .A(n377), .B(n376), .C(n375), .Z(n370) );
  COND2XL U2303 ( .A(n1697), .B(n1153), .C(n74), .D(n1152), .Z(n874) );
  COND2XL U2304 ( .A(n1586), .B(n1155), .C(n74), .D(n1154), .Z(n876) );
  CFA1X1 U2305 ( .A(n979), .B(n843), .CI(n1063), .CO(n571), .S(n572) );
  COND2X1 U2306 ( .A(n1119), .B(n97), .C(n95), .D(n1118), .Z(n843) );
  COND2X1 U2307 ( .A(n1747), .B(n1737), .C(n1814), .D(n1106), .Z(n832) );
  CIVXL U2308 ( .A(n1610), .Z(n337) );
  CFA1X1 U2309 ( .A(n933), .B(n803), .CI(n913), .CO(n573), .S(n574) );
  CFA1X1 U2310 ( .A(n908), .B(n830), .CI(n2116), .CO(n455), .S(n456) );
  CFA1X1 U2311 ( .A(n820), .B(n838), .CI(n1606), .CO(n459), .S(n460) );
  CIVXL U2312 ( .A(n2010), .Z(n2001) );
  CND2X1 U2313 ( .A(n349), .B(n2111), .Z(n2010) );
  CENXL U2314 ( .A(n2160), .B(n2168), .Z(n1121) );
  CENXL U2315 ( .A(n2155), .B(n2168), .Z(n1126) );
  CENXL U2316 ( .A(n2156), .B(n2168), .Z(n1125) );
  CENXL U2317 ( .A(n2154), .B(n2168), .Z(n1127) );
  CENXL U2318 ( .A(n2157), .B(n2168), .Z(n1124) );
  CENXL U2319 ( .A(n2152), .B(n2168), .Z(n1129) );
  CENXL U2320 ( .A(n1388), .B(n1863), .Z(n1166) );
  CENXL U2321 ( .A(n2161), .B(n1857), .Z(n1171) );
  CENXL U2322 ( .A(n2158), .B(n1857), .Z(n1174) );
  CENXL U2323 ( .A(n2159), .B(n1857), .Z(n1173) );
  CENXL U2324 ( .A(n1389), .B(n1863), .Z(n1167) );
  CENXL U2325 ( .A(n2160), .B(n1856), .Z(n1172) );
  CENXL U2326 ( .A(n2164), .B(n1856), .Z(n1168) );
  CENXL U2327 ( .A(n2163), .B(n1857), .Z(n1169) );
  CENXL U2328 ( .A(n2162), .B(n1863), .Z(n1170) );
  CENXL U2329 ( .A(n2157), .B(n1857), .Z(n1175) );
  CENXL U2330 ( .A(n2156), .B(n1856), .Z(n1176) );
  CENXL U2331 ( .A(n2153), .B(n1856), .Z(n1179) );
  CENXL U2332 ( .A(n2154), .B(n1857), .Z(n1178) );
  CENXL U2333 ( .A(n2152), .B(n1857), .Z(n1180) );
  CENXL U2334 ( .A(n2155), .B(n1856), .Z(n1177) );
  CENXL U2335 ( .A(n2151), .B(n1856), .Z(n1181) );
  COND2X1 U2336 ( .A(n1570), .B(n1183), .C(n66), .D(n1182), .Z(n903) );
  CND2X2 U2337 ( .A(n1989), .B(n1988), .Z(product[30]) );
  COND2X1 U2338 ( .A(n77), .B(n1438), .C(n74), .D(n1165), .Z(n806) );
  CFA1X1 U2339 ( .A(n1069), .B(n806), .CI(n961), .CO(n683), .S(n684) );
  CND2X2 U2340 ( .A(n2007), .B(n1970), .Z(n1971) );
  CND2X1 U2341 ( .A(n1969), .B(n235), .Z(n1972) );
  CND2X4 U2342 ( .A(n1971), .B(n1972), .Z(product[20]) );
  CIVX2 U2343 ( .A(n2007), .Z(n1969) );
  CIVX1 U2344 ( .A(n235), .Z(n1970) );
  COND1X1 U2345 ( .A(n286), .B(n282), .C(n283), .Z(n281) );
  CNR2XL U2346 ( .A(n1225), .B(n1815), .Z(n1977) );
  CENXL U2347 ( .A(n2151), .B(n2201), .Z(n1225) );
  CND2XL U2348 ( .A(n2025), .B(n260), .Z(n1979) );
  CND2X2 U2349 ( .A(n1978), .B(net179418), .Z(n1980) );
  CND2X2 U2350 ( .A(n1979), .B(n1980), .Z(product[16]) );
  CIVX2 U2351 ( .A(n2025), .Z(n1978) );
  CIVX2 U2352 ( .A(n260), .Z(net179418) );
  CAN2XL U2353 ( .A(n348), .B(n255), .Z(n2025) );
  COND2X1 U2354 ( .A(n97), .B(n1112), .C(n95), .D(n1111), .Z(n836) );
  CENX2 U2355 ( .A(n2138), .B(a[20]), .Z(n89) );
  COND2X1 U2356 ( .A(n69), .B(n1439), .C(n66), .D(n1184), .Z(n807) );
  CEO3X1 U2357 ( .A(n878), .B(n932), .C(n912), .Z(n552) );
  CIVDX3 U2358 ( .A(n3), .Z0(net179383), .Z1(net179382) );
  COND2X2 U2359 ( .A(n1109), .B(n1814), .C(n102), .D(n1434), .Z(n802) );
  CND2XL U2360 ( .A(n548), .B(n569), .Z(n2147) );
  CNR2X2 U2361 ( .A(n2034), .B(n2032), .Z(n254) );
  COND1X1 U2362 ( .A(n2097), .B(n262), .C(n263), .Z(n261) );
  CAN2XL U2363 ( .A(n335), .B(n163), .Z(n2016) );
  CIVXL U2364 ( .A(n230), .Z(n1992) );
  COND1X1 U2365 ( .A(n239), .B(n233), .C(n234), .Z(n232) );
  CIVXL U2366 ( .A(n131), .Z(n1995) );
  CEOXL U2367 ( .A(n2139), .B(n634), .Z(n626) );
  CNIVX3 U2368 ( .A(n1393), .Z(n2161) );
  CIVX2 U2369 ( .A(n182), .Z(n1999) );
  CIVXL U2370 ( .A(n184), .Z(n182) );
  CANR1X1 U2371 ( .A(n330), .B(n2023), .C(n327), .Z(n325) );
  CND2IXL U2372 ( .B(n205), .A(net178605), .Z(n196) );
  CND2IXL U2373 ( .B(n2110), .A(n2109), .Z(n136) );
  CND2XL U2374 ( .A(n345), .B(n239), .Z(n131) );
  CIVX1 U2375 ( .A(n2175), .Z(n2173) );
  CND2XL U2376 ( .A(n463), .B(n438), .Z(n2125) );
  CNIVX2 U2377 ( .A(n1392), .Z(n2162) );
  CNIVX2 U2378 ( .A(n1391), .Z(n2163) );
  CNIVX4 U2379 ( .A(n1397), .Z(n2157) );
  CND2XL U2380 ( .A(n1738), .B(n2001), .Z(n2002) );
  CND2XL U2381 ( .A(n2019), .B(n299), .Z(n141) );
  CND2XL U2382 ( .A(n2017), .B(n305), .Z(n142) );
  CND2IXL U2383 ( .B(n282), .A(n283), .Z(n138) );
  CENX1 U2384 ( .A(n2004), .B(n2005), .Z(product[24]) );
  CND2XL U2385 ( .A(net178605), .B(net179838), .Z(n2005) );
  CND2IXL U2386 ( .B(n307), .A(n308), .Z(n143) );
  CND2IXL U2387 ( .B(n315), .A(n316), .Z(n145) );
  CND2XL U2388 ( .A(n2022), .B(n313), .Z(n144) );
  CND2XL U2389 ( .A(n2023), .B(n329), .Z(n148) );
  CND2XL U2390 ( .A(n2021), .B(n321), .Z(n146) );
  CENXL U2391 ( .A(a[22]), .B(n93), .Z(n2006) );
  CENX1 U2392 ( .A(net178962), .B(n1612), .Z(product[22]) );
  CND2XL U2393 ( .A(n1590), .B(n184), .Z(n124) );
  CND2XL U2394 ( .A(n179), .B(n337), .Z(n123) );
  CEOX2 U2395 ( .A(n1928), .B(n1587), .Z(n1411) );
  CND2XL U2396 ( .A(n344), .B(n234), .Z(n2007) );
  CEOXL U2397 ( .A(n2132), .B(n551), .Z(n522) );
  CND2XL U2398 ( .A(n798), .B(n1053), .Z(n324) );
  CND2XL U2399 ( .A(n532), .B(n551), .Z(n2134) );
  CND2X2 U2400 ( .A(n2009), .B(n74), .Z(n77) );
  CIVX3 U2401 ( .A(n2198), .Z(n2193) );
  CENXL U2402 ( .A(n2161), .B(n2138), .Z(n1135) );
  COND2XL U2403 ( .A(n84), .B(n1140), .C(n82), .D(n1139), .Z(n862) );
  COND2X1 U2404 ( .A(n18), .B(n1338), .C(n1337), .D(n15), .Z(n1052) );
  CND2X2 U2405 ( .A(n353), .B(n2104), .Z(n139) );
  CNIVX2 U2406 ( .A(n1390), .Z(n2164) );
  CNIVX4 U2407 ( .A(n1400), .Z(n2154) );
  CENX1 U2408 ( .A(a[4]), .B(n2181), .Z(n2011) );
  CNIVX4 U2409 ( .A(n1402), .Z(n2152) );
  CNIVX4 U2410 ( .A(n1401), .Z(n2153) );
  CENX4 U2411 ( .A(n2178), .B(a[6]), .Z(net178746) );
  CANR1XL U2412 ( .A(n349), .B(n270), .C(n265), .Z(n263) );
  CND2XL U2413 ( .A(n269), .B(n349), .Z(n262) );
  CNIVX4 U2414 ( .A(n1398), .Z(n2156) );
  CIVX2 U2415 ( .A(n119), .Z(n2013) );
  CIVXL U2416 ( .A(n208), .Z(net178660) );
  COND1XL U2417 ( .A(n301), .B(n289), .C(n290), .Z(n288) );
  CENX1 U2418 ( .A(n141), .B(n300), .Z(product[9]) );
  CND2XL U2419 ( .A(n716), .B(n727), .Z(n272) );
  CND3XL U2420 ( .A(n2129), .B(n2130), .C(n2131), .Z(n551) );
  COND1XL U2421 ( .A(n196), .B(n1612), .C(n197), .Z(n195) );
  CANR1XL U2422 ( .A(net178605), .B(n208), .C(net180217), .Z(n197) );
  CENX1 U2423 ( .A(n144), .B(n314), .Z(product[6]) );
  CENX1 U2424 ( .A(n148), .B(n330), .Z(product[2]) );
  CENX1 U2425 ( .A(n146), .B(n322), .Z(product[4]) );
  CNR2X1 U2426 ( .A(n750), .B(n759), .Z(n285) );
  CEOXL U2427 ( .A(n325), .B(n147), .Z(product[3]) );
  CND2X1 U2428 ( .A(n361), .B(n324), .Z(n147) );
  COR2X1 U2429 ( .A(n776), .B(n781), .Z(n2017) );
  COR2X1 U2430 ( .A(n760), .B(n767), .Z(n2018) );
  CND2X1 U2431 ( .A(n768), .B(n775), .Z(n299) );
  CND2X1 U2432 ( .A(n776), .B(n781), .Z(n305) );
  CND2X1 U2433 ( .A(n760), .B(n767), .Z(n294) );
  CNR2X1 U2434 ( .A(n1553), .B(n739), .Z(n276) );
  COR2X1 U2435 ( .A(n768), .B(n775), .Z(n2019) );
  CND2X1 U2436 ( .A(n750), .B(n759), .Z(n286) );
  CND2XL U2437 ( .A(n728), .B(n739), .Z(n277) );
  COR2X1 U2438 ( .A(n380), .B(n407), .Z(n2020) );
  CEOXL U2439 ( .A(n636), .B(n632), .Z(n2139) );
  CNR2X1 U2440 ( .A(n792), .B(n795), .Z(n315) );
  CND3XL U2441 ( .A(n2140), .B(n2141), .C(n2142), .Z(n633) );
  CNR2X1 U2442 ( .A(n782), .B(n787), .Z(n307) );
  CNR2X1 U2443 ( .A(n798), .B(n1053), .Z(n323) );
  CND3XL U2444 ( .A(n2146), .B(n2147), .C(n2148), .Z(n541) );
  CND2X1 U2445 ( .A(n792), .B(n795), .Z(n316) );
  CND2X1 U2446 ( .A(n796), .B(n797), .Z(n321) );
  CND2X1 U2447 ( .A(n788), .B(n791), .Z(n313) );
  CND2X1 U2448 ( .A(n1084), .B(n1054), .Z(n329) );
  CND3XL U2449 ( .A(n2133), .B(n2134), .C(n2135), .Z(n521) );
  CND2X1 U2450 ( .A(n782), .B(n787), .Z(n308) );
  COR2X1 U2451 ( .A(n796), .B(n797), .Z(n2021) );
  COR2X1 U2452 ( .A(n788), .B(n791), .Z(n2022) );
  COR2X1 U2453 ( .A(n1084), .B(n1054), .Z(n2023) );
  CAN2XL U2454 ( .A(n1593), .B(n332), .Z(product[1]) );
  CENXL U2455 ( .A(n2151), .B(net183987), .Z(n1090) );
  CENXL U2456 ( .A(n2152), .B(net183987), .Z(n1089) );
  COR2X1 U2457 ( .A(n600), .B(n619), .Z(net178512) );
  CND3X1 U2458 ( .A(n2120), .B(n2121), .C(n2122), .Z(n437) );
  CND2X1 U2459 ( .A(n620), .B(n637), .Z(n234) );
  CND2X1 U2460 ( .A(n462), .B(n487), .Z(n179) );
  CND2X1 U2461 ( .A(n600), .B(n619), .Z(n229) );
  CND2X1 U2462 ( .A(n436), .B(n461), .Z(n170) );
  CENX1 U2463 ( .A(net33076), .B(n2172), .Z(n1339) );
  CENX1 U2464 ( .A(n2172), .B(n2159), .Z(n1329) );
  CENX1 U2465 ( .A(n2174), .B(n2158), .Z(n1330) );
  CENX1 U2466 ( .A(n2178), .B(n2158), .Z(n1299) );
  CENX1 U2467 ( .A(n2194), .B(n2161), .Z(n1240) );
  CENX1 U2468 ( .A(n2186), .B(n2164), .Z(n1264) );
  CENX1 U2469 ( .A(n2194), .B(n2164), .Z(n1237) );
  CENX1 U2470 ( .A(net179382), .B(net33422), .Z(n1371) );
  CENX1 U2471 ( .A(net179382), .B(n2151), .Z(n1370) );
  CENX1 U2472 ( .A(net179382), .B(n2153), .Z(n1368) );
  CENX1 U2473 ( .A(net179382), .B(n2152), .Z(n1369) );
  CENX1 U2474 ( .A(net179382), .B(n2155), .Z(n1366) );
  CENX1 U2475 ( .A(net179382), .B(n2157), .Z(n1364) );
  CENX1 U2476 ( .A(net179382), .B(n2158), .Z(n1363) );
  CENX1 U2477 ( .A(net179382), .B(n2160), .Z(n1361) );
  CENX1 U2478 ( .A(net179382), .B(n2156), .Z(n1365) );
  CENX1 U2479 ( .A(net179382), .B(n2159), .Z(n1362) );
  CENX1 U2480 ( .A(net179382), .B(n2154), .Z(n1367) );
  CENX1 U2481 ( .A(net32098), .B(n2164), .Z(n1357) );
  CENX2 U2482 ( .A(n2193), .B(a[10]), .Z(n50) );
  CENX1 U2483 ( .A(n2193), .B(n2157), .Z(n1244) );
  CENX1 U2484 ( .A(n2177), .B(n2153), .Z(n1304) );
  CENX1 U2485 ( .A(n2179), .B(n2161), .Z(n1296) );
  CENX1 U2486 ( .A(n2178), .B(n2159), .Z(n1298) );
  CENX1 U2487 ( .A(n2193), .B(n2158), .Z(n1243) );
  CENX1 U2488 ( .A(n2178), .B(n2157), .Z(n1300) );
  CENX1 U2489 ( .A(n2186), .B(n2163), .Z(n1265) );
  CENX1 U2490 ( .A(net33076), .B(net32098), .Z(n1372) );
  CENX1 U2491 ( .A(n2176), .B(n2155), .Z(n1302) );
  CENX1 U2492 ( .A(n2180), .B(n2156), .Z(n1301) );
  CENX1 U2493 ( .A(n2179), .B(n2154), .Z(n1303) );
  CENX1 U2494 ( .A(n2186), .B(n2162), .Z(n1266) );
  CNR2IXL U2495 ( .B(net33078), .A(n15), .Z(n1054) );
  CENX1 U2496 ( .A(n2173), .B(n2162), .Z(n1326) );
  CENX1 U2497 ( .A(n2179), .B(n2163), .Z(n1294) );
  CENX1 U2498 ( .A(n2180), .B(n2164), .Z(n1293) );
  CENX1 U2499 ( .A(n2194), .B(n2162), .Z(n1239) );
  CENX1 U2500 ( .A(n2194), .B(n2163), .Z(n1238) );
  CENX1 U2501 ( .A(n2185), .B(n2158), .Z(n1270) );
  CENX1 U2502 ( .A(n2170), .B(n2161), .Z(n1327) );
  CENX1 U2503 ( .A(n2170), .B(n2160), .Z(n1328) );
  CENX1 U2504 ( .A(n2151), .B(n2196), .Z(n1250) );
  CENX1 U2505 ( .A(n2185), .B(n2159), .Z(n1269) );
  CENX1 U2506 ( .A(n2173), .B(n2156), .Z(n1332) );
  CENX1 U2507 ( .A(n2170), .B(n2163), .Z(n1325) );
  CENX1 U2508 ( .A(n2194), .B(n2159), .Z(n1242) );
  CENX1 U2509 ( .A(n2177), .B(n2152), .Z(n1305) );
  CENX1 U2510 ( .A(n2192), .B(n2156), .Z(n1245) );
  CENX1 U2511 ( .A(n2179), .B(n2160), .Z(n1297) );
  CENX1 U2512 ( .A(n2183), .B(n2157), .Z(n1271) );
  CENX1 U2513 ( .A(n2173), .B(n2164), .Z(n1324) );
  CENX1 U2514 ( .A(n2179), .B(n2162), .Z(n1295) );
  CENX1 U2515 ( .A(n2194), .B(n2160), .Z(n1241) );
  CENXL U2516 ( .A(n2155), .B(n1933), .Z(n1113) );
  CENXL U2517 ( .A(n2160), .B(n2138), .Z(n1136) );
  CENX1 U2518 ( .A(net33076), .B(n2187), .Z(n1279) );
  CENX1 U2519 ( .A(n2177), .B(n2151), .Z(n1306) );
  CENX1 U2520 ( .A(n2172), .B(n2151), .Z(n1337) );
  CENX1 U2521 ( .A(n2177), .B(net33422), .Z(n1307) );
  CENX1 U2522 ( .A(n2172), .B(net33422), .Z(n1338) );
  CENX1 U2523 ( .A(n2184), .B(n2153), .Z(n1275) );
  CENX1 U2524 ( .A(n2184), .B(n2152), .Z(n1276) );
  CENX1 U2525 ( .A(n2183), .B(n2155), .Z(n1273) );
  CENX1 U2526 ( .A(n2184), .B(n2151), .Z(n1277) );
  CENX1 U2527 ( .A(n2184), .B(n2154), .Z(n1274) );
  CENX1 U2528 ( .A(n2172), .B(n2152), .Z(n1336) );
  CENX1 U2529 ( .A(n2152), .B(n2196), .Z(n1249) );
  CENX1 U2530 ( .A(n2173), .B(n2153), .Z(n1335) );
  CENX1 U2531 ( .A(n2185), .B(n2160), .Z(n1268) );
  CENX1 U2532 ( .A(n2170), .B(n2154), .Z(n1334) );
  CENX1 U2533 ( .A(n2183), .B(n2156), .Z(n1272) );
  CENX1 U2534 ( .A(n2192), .B(n2153), .Z(n1248) );
  CENX1 U2535 ( .A(n2183), .B(net33422), .Z(n1278) );
  CENX1 U2536 ( .A(n2192), .B(n2155), .Z(n1246) );
  CENX1 U2537 ( .A(n2192), .B(n2154), .Z(n1247) );
  CENX1 U2538 ( .A(n2185), .B(n2161), .Z(n1267) );
  CNR2X1 U2539 ( .A(n638), .B(n655), .Z(n238) );
  CENX1 U2540 ( .A(net33078), .B(n2181), .Z(n1308) );
  CND2X1 U2541 ( .A(n638), .B(n655), .Z(n239) );
  CND2X1 U2542 ( .A(n656), .B(n671), .Z(n245) );
  CIVX2 U2543 ( .A(net179383), .Z(net32098) );
  CND2X1 U2544 ( .A(n1592), .B(n151), .Z(n119) );
  CND2XL U2545 ( .A(n379), .B(n364), .Z(n151) );
  CNR2IXL U2546 ( .B(net33078), .A(n6), .Z(product[0]) );
  CND3X1 U2547 ( .A(net33752), .B(n2149), .C(net33754), .Z(n513) );
  CENX1 U2548 ( .A(n2027), .B(n493), .Z(n466) );
  CENX1 U2549 ( .A(n2073), .B(n2066), .Z(n2027) );
  CND3X1 U2550 ( .A(n2126), .B(n2127), .C(n2128), .Z(n465) );
  CND2X1 U2551 ( .A(n493), .B(n2066), .Z(n2126) );
  CND2X1 U2552 ( .A(n493), .B(n2073), .Z(n2127) );
  CENX1 U2553 ( .A(n2177), .B(b[27]), .Z(n1281) );
  CENX1 U2554 ( .A(n2174), .B(n1389), .Z(n1323) );
  CENX1 U2555 ( .A(n2170), .B(n1386), .Z(n1320) );
  CENX1 U2556 ( .A(n2187), .B(n1387), .Z(n1261) );
  CENX1 U2557 ( .A(net32098), .B(n1389), .Z(n1356) );
  CENX1 U2558 ( .A(net32098), .B(n1388), .Z(n1355) );
  CENX1 U2559 ( .A(net179382), .B(n1385), .Z(n1352) );
  CENX1 U2560 ( .A(net179382), .B(n1384), .Z(n1351) );
  CENX1 U2561 ( .A(net179382), .B(n1383), .Z(n1350) );
  CENX1 U2562 ( .A(net179382), .B(n1387), .Z(n1354) );
  CENX1 U2563 ( .A(net179382), .B(n1386), .Z(n1353) );
  CENX1 U2564 ( .A(net179382), .B(b[25]), .Z(n1347) );
  CENX1 U2565 ( .A(net179382), .B(b[29]), .Z(n1343) );
  CENX1 U2566 ( .A(net179382), .B(b[30]), .Z(n1342) );
  CENX1 U2567 ( .A(net179382), .B(b[24]), .Z(n1348) );
  CENX1 U2568 ( .A(net179382), .B(n1382), .Z(n1349) );
  CENX1 U2569 ( .A(net179382), .B(b[26]), .Z(n1346) );
  CENX1 U2570 ( .A(net179382), .B(b[28]), .Z(n1344) );
  CENX1 U2571 ( .A(net179382), .B(b[27]), .Z(n1345) );
  CENX1 U2572 ( .A(n2172), .B(n1388), .Z(n1322) );
  CENX1 U2573 ( .A(n2191), .B(n1385), .Z(n1232) );
  CENX1 U2574 ( .A(n2186), .B(n1389), .Z(n1263) );
  CENX1 U2575 ( .A(n2187), .B(n1388), .Z(n1262) );
  CENX1 U2576 ( .A(n2193), .B(n1382), .Z(n1229) );
  CENX1 U2577 ( .A(n2186), .B(b[25]), .Z(n1254) );
  CENX1 U2578 ( .A(net179382), .B(b[31]), .Z(n1341) );
  CENX1 U2579 ( .A(n2186), .B(n1383), .Z(n1257) );
  CENX1 U2580 ( .A(n2186), .B(n1382), .Z(n1256) );
  CENX1 U2581 ( .A(n2186), .B(b[24]), .Z(n1255) );
  CENX1 U2582 ( .A(n2172), .B(n1382), .Z(n1316) );
  CENX1 U2583 ( .A(n2180), .B(n1384), .Z(n1287) );
  CENX1 U2584 ( .A(n2194), .B(n1387), .Z(n1234) );
  CENX1 U2585 ( .A(n2180), .B(n1387), .Z(n1290) );
  CENX1 U2586 ( .A(n2194), .B(n1389), .Z(n1236) );
  CENX1 U2587 ( .A(n2173), .B(n1383), .Z(n1317) );
  CENX1 U2588 ( .A(n2180), .B(n1383), .Z(n1286) );
  CENX1 U2589 ( .A(n2172), .B(b[25]), .Z(n1314) );
  CENX1 U2590 ( .A(n2180), .B(n1382), .Z(n1285) );
  CENX1 U2591 ( .A(n2172), .B(b[26]), .Z(n1313) );
  CENX1 U2592 ( .A(n2180), .B(n1389), .Z(n1292) );
  CENX1 U2593 ( .A(n2176), .B(n1386), .Z(n1289) );
  CENX1 U2594 ( .A(n2176), .B(b[24]), .Z(n1284) );
  CENX1 U2595 ( .A(n2172), .B(b[27]), .Z(n1312) );
  CENX1 U2596 ( .A(n2180), .B(n1388), .Z(n1291) );
  CENX1 U2597 ( .A(n2180), .B(n1385), .Z(n1288) );
  CENX1 U2598 ( .A(n2183), .B(n1384), .Z(n1258) );
  CENX1 U2599 ( .A(n2191), .B(n1384), .Z(n1231) );
  CENX1 U2600 ( .A(n2191), .B(n1383), .Z(n1230) );
  CENX1 U2601 ( .A(n2176), .B(b[26]), .Z(n1282) );
  CENX1 U2602 ( .A(n2172), .B(b[28]), .Z(n1311) );
  CENX1 U2603 ( .A(n2176), .B(b[25]), .Z(n1283) );
  CENX1 U2604 ( .A(n2173), .B(b[29]), .Z(n1310) );
  CEO3X1 U2605 ( .A(n385), .B(n2028), .C(n2029), .Z(n365) );
  CEN3X2 U2606 ( .A(n2093), .B(n2095), .C(n2100), .Z(n2028) );
  CEN3X1 U2607 ( .A(n2101), .B(n387), .C(n368), .Z(n2029) );
  CNIVX4 U2608 ( .A(n1403), .Z(n2151) );
  CIVX2 U2609 ( .A(n39), .Z(n2198) );
  CNIVX4 U2610 ( .A(n1399), .Z(n2155) );
  CENX1 U2611 ( .A(n2175), .B(a[4]), .Z(n2030) );
  CIVX4 U2612 ( .A(n2030), .Z(n24) );
  CEOX2 U2613 ( .A(n30), .B(a[8]), .Z(n2031) );
  CIVX4 U2614 ( .A(n2031), .Z(n42) );
  CNIVX3 U2615 ( .A(n1394), .Z(n2160) );
  CNIVX4 U2616 ( .A(n1396), .Z(n2158) );
  CNIVX4 U2617 ( .A(n1395), .Z(n2159) );
  COND2XL U2618 ( .A(n1586), .B(n1150), .C(n74), .D(n1149), .Z(n871) );
  COND2XL U2619 ( .A(n1697), .B(n1151), .C(n74), .D(n1150), .Z(n872) );
  COND2XL U2620 ( .A(n1697), .B(n1158), .C(n74), .D(n1157), .Z(n879) );
  COND2XL U2621 ( .A(n1697), .B(n1152), .C(n74), .D(n1151), .Z(n873) );
  COND2XL U2622 ( .A(n1697), .B(n1154), .C(n74), .D(n1153), .Z(n875) );
  COND2XL U2623 ( .A(n77), .B(n1161), .C(n74), .D(n1160), .Z(n882) );
  COND2XL U2624 ( .A(n1697), .B(n1159), .C(n74), .D(n1158), .Z(n880) );
  CND2IXL U2625 ( .B(net33078), .A(n2168), .Z(n1133) );
  CENXL U2626 ( .A(n2159), .B(n2168), .Z(n1122) );
  CIVXL U2627 ( .A(n1672), .Z(n1438) );
  CIVXL U2628 ( .A(n890), .Z(n2115) );
  CIVX1 U2629 ( .A(n2115), .Z(n2116) );
  COND2XL U2630 ( .A(n91), .B(n1126), .C(n89), .D(n1125), .Z(n849) );
  CEOXL U2631 ( .A(n845), .B(n871), .Z(n378) );
  CNIVX1 U2632 ( .A(n927), .Z(n2118) );
  CFA1XL U2633 ( .A(n914), .B(n1064), .CI(n934), .CO(n593), .S(n594) );
  COND2XL U2634 ( .A(n36), .B(n1259), .C(n1258), .D(net178746), .Z(n975) );
  COND2XL U2635 ( .A(n36), .B(n1263), .C(n1262), .D(net178746), .Z(n979) );
  COND2XL U2636 ( .A(n36), .B(n1267), .C(n1266), .D(net178746), .Z(n983) );
  COND2XL U2637 ( .A(n36), .B(n1268), .C(n1267), .D(net178746), .Z(n984) );
  COND2XL U2638 ( .A(n36), .B(n1269), .C(n1268), .D(net178746), .Z(n985) );
  CNR2IXL U2639 ( .B(net33078), .A(net178746), .Z(n996) );
  COND2XL U2640 ( .A(n1279), .B(n36), .C(n1278), .D(net178746), .Z(n995) );
  COND2XL U2641 ( .A(n36), .B(n1277), .C(n1276), .D(net178746), .Z(n993) );
  COND2XL U2642 ( .A(n36), .B(n1275), .C(n1274), .D(net178746), .Z(n991) );
  COND2XL U2643 ( .A(n36), .B(n1273), .C(n1272), .D(net178746), .Z(n989) );
  COND2XL U2644 ( .A(n36), .B(n1272), .C(n1271), .D(net178746), .Z(n988) );
  COND2XL U2645 ( .A(n36), .B(n1255), .C(n1254), .D(net178746), .Z(n971) );
  COND2XL U2646 ( .A(n36), .B(n1266), .C(n1265), .D(net178746), .Z(n982) );
  CEO3X2 U2647 ( .A(n444), .B(n465), .C(n442), .Z(n438) );
  CEOX1 U2648 ( .A(n2119), .B(n438), .Z(n436) );
  CND2X1 U2649 ( .A(n444), .B(n465), .Z(n2120) );
  CND2X1 U2650 ( .A(n444), .B(n442), .Z(n2121) );
  CND2X1 U2651 ( .A(n465), .B(n442), .Z(n2122) );
  CND2XL U2652 ( .A(n440), .B(n463), .Z(n2123) );
  CND2X1 U2653 ( .A(n440), .B(n438), .Z(n2124) );
  CND2XL U2654 ( .A(n2066), .B(n2073), .Z(n2128) );
  COND2XL U2655 ( .A(n2117), .B(n1213), .C(n1212), .D(n1815), .Z(n931) );
  COND2XL U2656 ( .A(n53), .B(n1209), .C(n1208), .D(n1815), .Z(n927) );
  COND2XL U2657 ( .A(n53), .B(n1218), .C(n1217), .D(n1815), .Z(n936) );
  CIVXL U2658 ( .A(net179529), .Z(n208) );
  CFA1XL U2659 ( .A(n880), .B(n956), .CI(n896), .CO(n595), .S(n596) );
  CND2X1 U2660 ( .A(n380), .B(n407), .Z(n156) );
  CIVX1 U2661 ( .A(n156), .Z(n154) );
  CIVXL U2662 ( .A(n1986), .Z(n335) );
  CIVXL U2663 ( .A(n233), .Z(n344) );
  CIVXL U2664 ( .A(n1857), .Z(n1439) );
  CND2XL U2665 ( .A(n878), .B(n932), .Z(n2129) );
  CND2XL U2666 ( .A(n878), .B(n912), .Z(n2130) );
  CND2X1 U2667 ( .A(n932), .B(n912), .Z(n2131) );
  CND2X1 U2668 ( .A(n532), .B(n549), .Z(n2133) );
  CND2X1 U2669 ( .A(n549), .B(n551), .Z(n2135) );
  CNR2XL U2670 ( .A(n1586), .B(n1157), .Z(n2136) );
  CNR2XL U2671 ( .A(n74), .B(n1156), .Z(n2137) );
  COR2X1 U2672 ( .A(n2136), .B(n2137), .Z(n878) );
  CIVX2 U2673 ( .A(n2175), .Z(n2171) );
  CIVX1 U2674 ( .A(n2175), .Z(n2170) );
  CIVX2 U2675 ( .A(n2175), .Z(n2172) );
  COND2XL U2676 ( .A(n84), .B(n1137), .C(n82), .D(n1136), .Z(n859) );
  COND2XL U2677 ( .A(n1147), .B(n84), .C(n82), .D(n1146), .Z(n869) );
  COND2XL U2678 ( .A(n84), .B(n1135), .C(n82), .D(n1134), .Z(n857) );
  CNR2X1 U2679 ( .A(n580), .B(n599), .Z(n216) );
  CNR2X1 U2680 ( .A(n233), .B(n238), .Z(n231) );
  CFA1XL U2681 ( .A(n918), .B(n1068), .CI(n960), .CO(n667), .S(n668) );
  CFA1X1 U2682 ( .A(n1584), .B(n1060), .CI(n976), .CO(n503), .S(n504) );
  COND2XL U2683 ( .A(n9), .B(net179383), .C(n6), .D(n1373), .Z(n814) );
  CND2X1 U2684 ( .A(n1085), .B(n814), .Z(n332) );
  CENX1 U2685 ( .A(net32098), .B(n2161), .Z(n1360) );
  CENX1 U2686 ( .A(net32098), .B(n2162), .Z(n1359) );
  CENX1 U2687 ( .A(net32098), .B(n2163), .Z(n1358) );
  CND2IXL U2688 ( .B(net33078), .A(net32098), .Z(n1373) );
  CENXL U2689 ( .A(n1696), .B(n1387), .Z(n1186) );
  CENXL U2690 ( .A(n2203), .B(n1388), .Z(n1187) );
  CIVX1 U2691 ( .A(n2205), .Z(n2204) );
  COND2XL U2692 ( .A(n27), .B(n1282), .C(n1281), .D(n24), .Z(n997) );
  COND2XL U2693 ( .A(n27), .B(n1283), .C(n1282), .D(n24), .Z(n998) );
  COND2XL U2694 ( .A(n27), .B(n1304), .C(n1303), .D(n24), .Z(n1019) );
  COND2XL U2695 ( .A(n27), .B(n1301), .C(n1300), .D(n24), .Z(n1016) );
  COND2XL U2696 ( .A(n1308), .B(n27), .C(n1307), .D(n24), .Z(n1023) );
  COND2XL U2697 ( .A(n27), .B(n1289), .C(n1288), .D(n24), .Z(n1004) );
  COND2XL U2698 ( .A(n27), .B(n2182), .C(n24), .D(n1309), .Z(n812) );
  COND2XL U2699 ( .A(n27), .B(n1298), .C(n1297), .D(n24), .Z(n1013) );
  COND2XL U2700 ( .A(n27), .B(n1296), .C(n1295), .D(n24), .Z(n1011) );
  COND2XL U2701 ( .A(n27), .B(n1284), .C(n1283), .D(n24), .Z(n999) );
  COND2XL U2702 ( .A(n27), .B(n1292), .C(n1291), .D(n24), .Z(n1007) );
  COND2XL U2703 ( .A(n27), .B(n1307), .C(n1306), .D(n24), .Z(n1022) );
  CND2XL U2704 ( .A(n2018), .B(n2019), .Z(n289) );
  CND2IXL U2705 ( .B(net33078), .A(n1672), .Z(n1165) );
  COND2X1 U2706 ( .A(n2117), .B(n1223), .C(n1222), .D(n1816), .Z(n941) );
  CND2IXL U2707 ( .B(net33078), .A(n1857), .Z(n1184) );
  COND2XL U2708 ( .A(n91), .B(n1122), .C(n89), .D(n1121), .Z(n845) );
  CHA1XL U2709 ( .A(n865), .B(n895), .CO(n577), .S(n578) );
  COND2XL U2710 ( .A(n77), .B(n1162), .C(n74), .D(n1161), .Z(n883) );
  COND2XL U2711 ( .A(n84), .B(n1143), .C(n82), .D(n1142), .Z(n865) );
  COND2XL U2712 ( .A(n84), .B(n1142), .C(n82), .D(n1141), .Z(n864) );
  CIVX1 U2713 ( .A(n2189), .Z(n2184) );
  CFA1XL U2714 ( .A(n940), .B(n1070), .CI(n1012), .CO(n697), .S(n698) );
  CIVX2 U2715 ( .A(n2190), .Z(n2185) );
  CIVX1 U2716 ( .A(n2190), .Z(n2186) );
  COND2XL U2717 ( .A(n1585), .B(n1167), .C(n1166), .D(n1596), .Z(n887) );
  COND2XL U2718 ( .A(n1585), .B(n1169), .C(n66), .D(n1168), .Z(n889) );
  COND2XL U2719 ( .A(n1585), .B(n1168), .C(n1167), .D(n1596), .Z(n888) );
  COND2XL U2720 ( .A(n1932), .B(n1181), .C(n66), .D(n1180), .Z(n901) );
  COND2XL U2721 ( .A(n1585), .B(n1174), .C(n1596), .D(n1173), .Z(n894) );
  COND2XL U2722 ( .A(n1585), .B(n1176), .C(n1596), .D(n1175), .Z(n896) );
  COND2XL U2723 ( .A(n1585), .B(n1170), .C(n1596), .D(n1169), .Z(n890) );
  COND2XL U2724 ( .A(n1585), .B(n1171), .C(n1596), .D(n1170), .Z(n891) );
  COND2XL U2725 ( .A(n1585), .B(n1173), .C(n66), .D(n1172), .Z(n893) );
  COND2XL U2726 ( .A(n1585), .B(n1175), .C(n1596), .D(n1174), .Z(n895) );
  COND2XL U2727 ( .A(n1932), .B(n1178), .C(n66), .D(n1177), .Z(n898) );
  CEO3XL U2728 ( .A(n898), .B(n1036), .C(n916), .Z(n634) );
  CND2XL U2729 ( .A(n898), .B(n1036), .Z(n2140) );
  CND2XL U2730 ( .A(n1036), .B(n916), .Z(n2142) );
  CND2X1 U2731 ( .A(n636), .B(n632), .Z(n2143) );
  CND2X1 U2732 ( .A(n636), .B(n634), .Z(n2144) );
  CND2X1 U2733 ( .A(n632), .B(n634), .Z(n2145) );
  CIVX1 U2734 ( .A(n2182), .Z(n2181) );
  CIVX2 U2735 ( .A(n2198), .Z(n2192) );
  COND1XL U2736 ( .A(n260), .B(n247), .C(n248), .Z(n246) );
  CND2XL U2737 ( .A(n514), .B(n516), .Z(n2150) );
  CIVX2 U2738 ( .A(n30), .Z(n2190) );
  COND2XL U2739 ( .A(n18), .B(n1322), .C(n1321), .D(n15), .Z(n1036) );
  CENX1 U2740 ( .A(n2191), .B(n1386), .Z(n1233) );
  CIVX2 U2741 ( .A(n2197), .Z(n2191) );
  COND2XL U2742 ( .A(net184278), .B(n1186), .C(n1185), .D(net180674), .Z(n905)
         );
  COND2XL U2743 ( .A(net184278), .B(n1187), .C(n1186), .D(net180674), .Z(n906)
         );
  COND2XL U2744 ( .A(net184278), .B(n1190), .C(n1189), .D(net180674), .Z(n909)
         );
  COND2XL U2745 ( .A(net184278), .B(n1189), .C(n1188), .D(net180674), .Z(n908)
         );
  COND2XL U2746 ( .A(n61), .B(n1201), .C(n58), .D(n1200), .Z(n920) );
  COND2XL U2747 ( .A(n61), .B(n1200), .C(n58), .D(n1199), .Z(n919) );
  COND2XL U2748 ( .A(n1599), .B(n1195), .C(n1194), .D(net180674), .Z(n914) );
  COND2XL U2749 ( .A(net184278), .B(n1194), .C(n1193), .D(net180674), .Z(n913)
         );
  COND2XL U2750 ( .A(n1599), .B(n1197), .C(net180674), .D(n1196), .Z(n916) );
  COND2XL U2751 ( .A(net184278), .B(n1191), .C(n1190), .D(net180674), .Z(n910)
         );
  COND2XL U2752 ( .A(n61), .B(n1198), .C(net180674), .D(n1197), .Z(n917) );
  COND2XL U2753 ( .A(net184278), .B(n1193), .C(n1192), .D(net180674), .Z(n912)
         );
  CENX1 U2754 ( .A(n2172), .B(n1385), .Z(n1319) );
  COND2X1 U2755 ( .A(n18), .B(n1315), .C(n1314), .D(n15), .Z(n1029) );
  CENX1 U2756 ( .A(n2183), .B(n1385), .Z(n1259) );
  CFA1XL U2757 ( .A(n915), .B(n1065), .CI(n935), .CO(n613), .S(n614) );
  CIVX1 U2758 ( .A(n2182), .Z(n2179) );
  CIVX1 U2759 ( .A(n2182), .Z(n2176) );
  CIVX1 U2760 ( .A(n2182), .Z(n2180) );
  CIVX1 U2761 ( .A(n2182), .Z(n2177) );
  COND2XL U2762 ( .A(n18), .B(n1311), .C(n1310), .D(n15), .Z(n1025) );
  COND2XL U2763 ( .A(n18), .B(n1312), .C(n1311), .D(n15), .Z(n1026) );
  COND2XL U2764 ( .A(n1339), .B(n18), .C(n1338), .D(n15), .Z(n1053) );
  COND2XL U2765 ( .A(n18), .B(n1337), .C(n1336), .D(n15), .Z(n1051) );
  COND2XL U2766 ( .A(n18), .B(n1335), .C(n1334), .D(n15), .Z(n1049) );
  COND2XL U2767 ( .A(n18), .B(n2175), .C(n15), .D(n1340), .Z(n813) );
  COND2XL U2768 ( .A(n18), .B(n1325), .C(n1324), .D(n15), .Z(n1039) );
  COND2XL U2769 ( .A(n18), .B(n1332), .C(n1331), .D(n15), .Z(n1046) );
  COND2XL U2770 ( .A(n18), .B(n1336), .C(n1335), .D(n15), .Z(n1050) );
  COND2XL U2771 ( .A(n18), .B(n1319), .C(n1318), .D(n15), .Z(n1033) );
  COND2XL U2772 ( .A(n36), .B(n2188), .C(net178746), .D(n1280), .Z(n811) );
  CND2IXL U2773 ( .B(net33078), .A(n2183), .Z(n1280) );
  CENX1 U2774 ( .A(n2186), .B(n1386), .Z(n1260) );
  COND2XL U2775 ( .A(n44), .B(n1230), .C(n1229), .D(n42), .Z(n947) );
  COND2XL U2776 ( .A(n44), .B(n1232), .C(n1231), .D(n42), .Z(n949) );
  COND2XL U2777 ( .A(n44), .B(n1231), .C(n1230), .D(n42), .Z(n948) );
  COND2XL U2778 ( .A(n44), .B(n2197), .C(n42), .D(n1253), .Z(n810) );
  COND2XL U2779 ( .A(n1252), .B(n44), .C(n1251), .D(n42), .Z(n969) );
  COND2XL U2780 ( .A(n44), .B(n1247), .C(n1246), .D(n42), .Z(n964) );
  COND2XL U2781 ( .A(n44), .B(n1246), .C(n1245), .D(n42), .Z(n963) );
  COND2XL U2782 ( .A(n44), .B(n1248), .C(n1247), .D(n42), .Z(n965) );
  COND2XL U2783 ( .A(n44), .B(n1242), .C(n1241), .D(n42), .Z(n959) );
  COND2XL U2784 ( .A(n44), .B(n1244), .C(n1243), .D(n42), .Z(n961) );
  CIVX1 U2785 ( .A(n2199), .Z(n2194) );
  CEOXL U2786 ( .A(n1959), .B(n143), .Z(product[7]) );
  CEOXL U2787 ( .A(n317), .B(n145), .Z(product[5]) );
  COND2XL U2788 ( .A(n2117), .B(n1207), .C(n1206), .D(n1815), .Z(n925) );
  COND2XL U2789 ( .A(n2117), .B(n1208), .C(n1207), .D(n1815), .Z(n926) );
  CNR2IXL U2790 ( .B(net33078), .A(n50), .Z(n946) );
  COND2XL U2791 ( .A(n2117), .B(n1210), .C(n1209), .D(n1815), .Z(n928) );
  COND2XL U2792 ( .A(n2117), .B(n1211), .C(n1210), .D(n1816), .Z(n929) );
  COND2XL U2793 ( .A(n2117), .B(n1220), .C(n1219), .D(n1815), .Z(n938) );
  COND2XL U2794 ( .A(n2117), .B(n1221), .C(n1220), .D(n1815), .Z(n939) );
  COND2XL U2795 ( .A(n2117), .B(n1215), .C(n1214), .D(n1816), .Z(n933) );
  COND2XL U2796 ( .A(n2117), .B(n1216), .C(n1215), .D(n1816), .Z(n934) );
  COND2XL U2797 ( .A(n2117), .B(n1668), .C(n1816), .D(n1224), .Z(n943) );
  COND2XL U2798 ( .A(n53), .B(n1222), .C(n1221), .D(n1815), .Z(n940) );
  COND2XL U2799 ( .A(n2117), .B(n1214), .C(n1213), .D(n1816), .Z(n932) );
  CND2X4 U2800 ( .A(n1421), .B(n6), .Z(n9) );
  CENX4 U2801 ( .A(n3), .B(a[2]), .Z(n15) );
  CND2X4 U2802 ( .A(n1420), .B(n15), .Z(n18) );
  CND2X4 U2803 ( .A(n1418), .B(net178746), .Z(n36) );
  CIVXL U2804 ( .A(n2175), .Z(n2174) );
  CIVXL U2805 ( .A(n30), .Z(n2188) );
  CIVXL U2806 ( .A(n2199), .Z(n2196) );
  CIVXL U2807 ( .A(n39), .Z(n2197) );
  CIVX2 U2808 ( .A(n323), .Z(n361) );
  CIVX2 U2809 ( .A(n2105), .Z(n353) );
  CIVX2 U2810 ( .A(n332), .Z(n330) );
  CIVX2 U2811 ( .A(n329), .Z(n327) );
  CIVX2 U2812 ( .A(n321), .Z(n319) );
  CIVX2 U2813 ( .A(n305), .Z(n303) );
  CIVX2 U2814 ( .A(n299), .Z(n297) );
  CIVX2 U2815 ( .A(n294), .Z(n292) );
  CIVX2 U2816 ( .A(n2112), .Z(n349) );
  CIVX2 U2817 ( .A(n254), .Z(n348) );
  CIVX2 U2818 ( .A(n239), .Z(n237) );
  CIVX2 U2819 ( .A(n238), .Z(n345) );
endmodule


module calc_DW02_mult_2_stage_1 ( A, B, TC, CLK, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC, CLK;
  wire   n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         \A_extended[32] , \B_extended[32] ;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33;
  assign \A_extended[32]  = A[31];
  assign \B_extended[32]  = B[31];

  calc_DW_mult_tc_22 mult_96 ( .a({\A_extended[32] , \A_extended[32] , A[30:0]}), .b({\B_extended[32] , \B_extended[32] , B[30:0]}), .product({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, PRODUCT[31:11], 
        n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26}), 
        .i_retiming_group_0_clk(CLK) );
  CFD1QX1 clk_r_REG207_S1 ( .D(n17), .CP(CLK), .Q(PRODUCT[9]) );
  CFD1QX1 clk_r_REG249_S1 ( .D(n18), .CP(CLK), .Q(PRODUCT[8]) );
  CFD1QX1 clk_r_REG261_S1 ( .D(n20), .CP(CLK), .Q(PRODUCT[6]) );
  CFD1QX1 clk_r_REG268_S1 ( .D(n22), .CP(CLK), .Q(PRODUCT[4]) );
  CFD1QX1 clk_r_REG273_S1 ( .D(n24), .CP(CLK), .Q(PRODUCT[2]) );
  CFD1QX1 clk_r_REG279_S1 ( .D(n25), .CP(CLK), .Q(PRODUCT[1]) );
  CFD1QX1 clk_r_REG281_S1 ( .D(n26), .CP(CLK), .Q(PRODUCT[0]) );
  CFD1QX2 clk_r_REG208_S1 ( .D(n16), .CP(CLK), .Q(PRODUCT[10]) );
  CFD1QX4 clk_r_REG258_S1 ( .D(n19), .CP(CLK), .Q(PRODUCT[7]) );
  CFD1QX4 clk_r_REG267_S1 ( .D(n21), .CP(CLK), .Q(PRODUCT[5]) );
  CFD1QX4 clk_r_REG271_S1 ( .D(n23), .CP(CLK), .Q(PRODUCT[3]) );
endmodule


module calc_DW_mult_tc_25 ( a, b, product, i_retiming_group_0_clk );
  input [32:0] a;
  input [32:0] b;
  output [65:0] product;
  input i_retiming_group_0_clk;
  wire   n6, n12, n18, n21, n24, n27, n30, n33, n36, n39, n42, n44, n48, n50,
         n53, n55, n58, n61, n63, n66, n69, n71, n74, n77, n79, n84, n86, n89,
         n91, n93, n95, n97, n99, n100, n102, n104, n105, n107, n109, n110,
         n112, n113, n114, n115, n116, n122, n124, n126, n127, n129, n131,
         n132, n133, n136, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n150, n152, n154, n156, n171, n172, n173, n176,
         n179, n187, n188, n192, n193, n204, n206, n213, n214, n216, n225,
         n233, n234, n238, n239, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n254, n256, n257, n258, n259, n261, n264,
         n265, n266, n267, n269, n271, n272, n273, n274, n275, n276, n279,
         n280, n281, n283, n284, n285, n286, n287, n289, n290, n291, n292,
         n293, n294, n296, n298, n299, n301, n303, n304, n305, n307, n309,
         n310, n311, n312, n313, n315, n317, n318, n319, n320, n321, n323,
         n325, n326, n327, n328, n329, n331, n333, n335, n347, n348, n349,
         n350, n352, n355, n357, n363, n365, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1410,
         n1411, n1412, n1413, n1414, n1417, n1419, n1421, n1422, n1423, n1424,
         n1435, n1436, n1437, net171532, net171533, net171534, net171535,
         net171536, net171537, net171538, net171539, net171540, net178944,
         net178945, net179451, net179450, net179577, net179704, net179703,
         net180090, net180181, net180264, net180393, net180512, net180533,
         net182652, net182753, net178510, n160, n158, net181713, net178506,
         n340, n168, n167, n166, n165, n163, net179550, n343, n342, n182, n181,
         n125, n226, net179908, net179873, net178516, net178515, n562, n561,
         n346, n228, n222, n215, n212, n210, n203, n201, n199, n198, n197,
         n196, net180047, net180046, net180045, net180044, net179917, n341,
         n195, n194, n184, n180, n175, n174, n170, n169, net179871, net179596,
         n604, n603, n584, n583, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876;
  assign n12 = a[3];
  assign n21 = a[5];
  assign n30 = a[7];
  assign n39 = a[9];
  assign n48 = a[11];
  assign n55 = a[13];
  assign n63 = a[15];
  assign n71 = a[17];
  assign n79 = a[19];
  assign n86 = a[21];
  assign n93 = a[23];
  assign n99 = a[25];
  assign n104 = a[27];
  assign n109 = a[29];
  assign n113 = a[32];
  assign n116 = b[0];
  assign n1386 = b[23];
  assign n1387 = b[22];
  assign n1388 = b[21];
  assign n1389 = b[20];
  assign n1390 = b[19];
  assign n1391 = b[18];
  assign n1392 = b[17];
  assign n1393 = b[16];
  assign n1394 = b[15];
  assign n1395 = b[14];
  assign n1396 = b[13];
  assign n1397 = b[12];
  assign n1398 = b[11];
  assign n1399 = b[10];
  assign n1400 = b[9];
  assign n1401 = b[8];
  assign n1402 = b[7];
  assign n1403 = b[6];
  assign n1404 = b[5];
  assign n1405 = b[4];
  assign n1406 = b[3];
  assign n1407 = b[2];
  assign n1408 = b[1];
  assign n1774 = i_retiming_group_0_clk;

  CNR2X2 U138 ( .A(n466), .B(n491), .Z(n176) );
  CNR2X2 U235 ( .A(n1723), .B(n1722), .Z(n248) );
  CND2X2 U295 ( .A(n357), .B(n1760), .Z(n139) );
  CEO3X2 U375 ( .A(n1750), .B(n1755), .C(n1752), .Z(n368) );
  CEO3X2 U376 ( .A(n389), .B(n371), .C(n370), .Z(n369) );
  CEO3X2 U377 ( .A(n373), .B(n391), .C(n372), .Z(n370) );
  CEO3X2 U378 ( .A(n375), .B(n374), .C(n393), .Z(n371) );
  CEO3X2 U379 ( .A(n397), .B(n376), .C(n395), .Z(n372) );
  CEO3X2 U382 ( .A(n405), .B(n401), .C(n381), .Z(n375) );
  CEO3X2 U383 ( .A(n409), .B(n382), .C(n407), .Z(n376) );
  CEO3X2 U388 ( .A(n821), .B(n831), .C(n839), .Z(n381) );
  CFA1X1 U390 ( .A(n1749), .B(n1751), .CI(n1748), .CO(n383), .S(n384) );
  CFA1X1 U391 ( .A(n392), .B(n415), .CI(n390), .CO(n385), .S(n386) );
  CFA1X1 U392 ( .A(n394), .B(n417), .CI(n419), .CO(n387), .S(n388) );
  CFA1X1 U393 ( .A(n398), .B(n396), .CI(n421), .CO(n389), .S(n390) );
  CFA1X1 U394 ( .A(n425), .B(n400), .CI(n423), .CO(n391), .S(n392) );
  CFA1X1 U395 ( .A(n427), .B(n402), .CI(n404), .CO(n393), .S(n394) );
  CFA1X1 U396 ( .A(n410), .B(n406), .CI(n408), .CO(n395), .S(n396) );
  CFA1X1 U397 ( .A(n433), .B(n429), .CI(n431), .CO(n397), .S(n398) );
  CFA1X1 U398 ( .A(n930), .B(n435), .CI(n437), .CO(n399), .S(n400) );
  CFA1X1 U399 ( .A(n910), .B(n1030), .CI(n952), .CO(n401), .S(n402) );
  CFA1X1 U400 ( .A(n892), .B(n1060), .CI(n976), .CO(n403), .S(n404) );
  CFA1X1 U402 ( .A(n876), .B(n832), .CI(n840), .CO(n407), .S(n408) );
  CFA1X1 U403 ( .A(n820), .B(n826), .CI(n822), .CO(n409), .S(n410) );
  CFA1X1 U404 ( .A(n1746), .B(n1747), .CI(n1745), .CO(n411), .S(n412) );
  CFA1X1 U405 ( .A(n420), .B(n443), .CI(n418), .CO(n413), .S(n414) );
  CFA1X1 U406 ( .A(n422), .B(n445), .CI(n447), .CO(n415), .S(n416) );
  CFA1X1 U407 ( .A(n426), .B(n424), .CI(n449), .CO(n417), .S(n418) );
  CFA1X1 U408 ( .A(n428), .B(n451), .CI(n453), .CO(n419), .S(n420) );
  CFA1X1 U410 ( .A(n457), .B(n436), .CI(n455), .CO(n423), .S(n424) );
  CFA1X1 U411 ( .A(n463), .B(n459), .CI(n461), .CO(n425), .S(n426) );
  CFA1X1 U412 ( .A(n953), .B(n438), .CI(n977), .CO(n427), .S(n428) );
  CFA1X1 U413 ( .A(n931), .B(n1031), .CI(n1003), .CO(n429), .S(n430) );
  CFA1X1 U415 ( .A(n823), .B(n911), .CI(n851), .CO(n433), .S(n434) );
  CFA1X1 U416 ( .A(n877), .B(n1577), .CI(n841), .CO(n435), .S(n436) );
  CHA1X1 U417 ( .A(n804), .B(n827), .CO(n437), .S(n438) );
  CFA1X1 U418 ( .A(n1743), .B(n1744), .CI(n1742), .CO(n439), .S(n440) );
  CFA1X1 U419 ( .A(n448), .B(n469), .CI(n446), .CO(n441), .S(n442) );
  CFA1X1 U420 ( .A(n450), .B(n471), .CI(n473), .CO(n443), .S(n444) );
  CFA1X1 U422 ( .A(n458), .B(n477), .CI(n479), .CO(n447), .S(n448) );
  CFA1X1 U424 ( .A(n481), .B(n464), .CI(n483), .CO(n451), .S(n452) );
  CFA1X1 U427 ( .A(n878), .B(n1032), .CI(n954), .CO(n457), .S(n458) );
  CFA1X1 U430 ( .A(n824), .B(n834), .CI(n828), .CO(n463), .S(n464) );
  CFA1X1 U431 ( .A(n1740), .B(n1741), .CI(n1739), .CO(n465), .S(n466) );
  CFA1X1 U432 ( .A(n474), .B(n495), .CI(n472), .CO(n467), .S(n468) );
  CFA1X1 U433 ( .A(n499), .B(n497), .CI(n476), .CO(n469), .S(n470) );
  CFA1X1 U434 ( .A(n480), .B(n478), .CI(n501), .CO(n471), .S(n472) );
  CFA1X1 U435 ( .A(n484), .B(n503), .CI(n482), .CO(n473), .S(n474) );
  CFA1X1 U437 ( .A(n511), .B(n507), .CI(n509), .CO(n477), .S(n478) );
  CFA1X1 U438 ( .A(n933), .B(n513), .CI(n490), .CO(n479), .S(n480) );
  CFA1X1 U439 ( .A(n1033), .B(n955), .CI(n913), .CO(n481), .S(n482) );
  CFA1X1 U440 ( .A(n1063), .B(n895), .CI(n979), .CO(n483), .S(n484) );
  CFA1X1 U441 ( .A(n865), .B(n1005), .CI(n853), .CO(n485), .S(n486) );
  CFA1X1 U442 ( .A(n879), .B(n829), .CI(n835), .CO(n487), .S(n488) );
  CHA1X1 U443 ( .A(n843), .B(n805), .CO(n489), .S(n490) );
  CFA1X1 U444 ( .A(n1737), .B(n1738), .CI(n1736), .CO(n491), .S(n492) );
  CFA1X1 U445 ( .A(n521), .B(n519), .CI(n498), .CO(n493), .S(n494) );
  CFA1X1 U446 ( .A(n523), .B(n500), .CI(n502), .CO(n495), .S(n496) );
  CFA1X1 U447 ( .A(n527), .B(n504), .CI(n525), .CO(n497), .S(n498) );
  CFA1X1 U448 ( .A(n510), .B(n506), .CI(n508), .CO(n499), .S(n500) );
  CFA1X1 U449 ( .A(n531), .B(n512), .CI(n514), .CO(n501), .S(n502) );
  CFA1X1 U450 ( .A(n535), .B(n529), .CI(n533), .CO(n503), .S(n504) );
  CFA1X1 U452 ( .A(n896), .B(n1034), .CI(n980), .CO(n507), .S(n508) );
  CFA1X1 U453 ( .A(n866), .B(n1064), .CI(n914), .CO(n509), .S(n510) );
  CFA1X1 U455 ( .A(n1778), .B(n844), .CI(n836), .CO(n513), .S(n514) );
  CFA1X1 U456 ( .A(n1734), .B(n1735), .CI(n1733), .CO(n515), .S(n516) );
  CFA1X1 U457 ( .A(n545), .B(n543), .CI(n522), .CO(n517), .S(n518) );
  CFA1X1 U458 ( .A(n526), .B(n547), .CI(n524), .CO(n519), .S(n520) );
  CFA1X1 U459 ( .A(n551), .B(n528), .CI(n549), .CO(n521), .S(n522) );
  CFA1X1 U460 ( .A(n534), .B(n530), .CI(n532), .CO(n523), .S(n524) );
  CFA1X1 U461 ( .A(n553), .B(n536), .CI(n555), .CO(n525), .S(n526) );
  CFA1X1 U463 ( .A(n897), .B(n1007), .CI(n981), .CO(n529), .S(n530) );
  CFA1X1 U464 ( .A(n881), .B(n1035), .CI(n957), .CO(n531), .S(n532) );
  CFA1X1 U465 ( .A(n1065), .B(n867), .CI(n915), .CO(n533), .S(n534) );
  CFA1X1 U466 ( .A(n837), .B(n935), .CI(n845), .CO(n535), .S(n536) );
  CHA1X1 U467 ( .A(n806), .B(n855), .CO(n537), .S(n538) );
  CFA1X1 U469 ( .A(n567), .B(n565), .CI(n546), .CO(n541), .S(n542) );
  CFA1X1 U470 ( .A(n569), .B(n548), .CI(n550), .CO(n543), .S(n544) );
  CFA1X1 U471 ( .A(n556), .B(n552), .CI(n571), .CO(n545), .S(n546) );
  CFA1X1 U472 ( .A(n558), .B(n573), .CI(n554), .CO(n547), .S(n548) );
  CFA1X1 U473 ( .A(n577), .B(n560), .CI(n575), .CO(n549), .S(n550) );
  CFA1X1 U474 ( .A(n936), .B(n579), .CI(n581), .CO(n551), .S(n552) );
  CFA1X1 U475 ( .A(n898), .B(n1008), .CI(n982), .CO(n553), .S(n554) );
  CFA1X1 U476 ( .A(n882), .B(n1036), .CI(n958), .CO(n555), .S(n556) );
  CFA1X1 U478 ( .A(n838), .B(n856), .CI(n846), .CO(n559), .S(n560) );
  CFA1X1 U480 ( .A(n570), .B(n587), .CI(n568), .CO(n563), .S(n564) );
  CFA1X1 U481 ( .A(n591), .B(n589), .CI(n572), .CO(n565), .S(n566) );
  CFA1X1 U482 ( .A(n576), .B(n574), .CI(n593), .CO(n567), .S(n568) );
  CFA1X1 U483 ( .A(n595), .B(n578), .CI(n580), .CO(n569), .S(n570) );
  CFA1X1 U484 ( .A(n601), .B(n597), .CI(n599), .CO(n571), .S(n572) );
  CFA1X1 U485 ( .A(n937), .B(n582), .CI(n959), .CO(n573), .S(n574) );
  CFA1X1 U487 ( .A(n857), .B(n983), .CI(n899), .CO(n577), .S(n578) );
  CFA1X1 U488 ( .A(n847), .B(n1009), .CI(n883), .CO(n579), .S(n580) );
  CFA1X1 U491 ( .A(n592), .B(n607), .CI(n590), .CO(n585), .S(n586) );
  CFA1X1 U492 ( .A(n611), .B(n609), .CI(n594), .CO(n587), .S(n588) );
  CFA1X1 U493 ( .A(n598), .B(n613), .CI(n596), .CO(n589), .S(n590) );
  CFA1X1 U494 ( .A(n617), .B(n600), .CI(n602), .CO(n591), .S(n592) );
  CFA1X1 U495 ( .A(n621), .B(n615), .CI(n619), .CO(n593), .S(n594) );
  CFA1X1 U497 ( .A(n1601), .B(n1589), .CI(n1010), .CO(n597), .S(n598) );
  CFA1X1 U499 ( .A(n848), .B(n870), .CI(n858), .CO(n601), .S(n602) );
  CFA1X1 U501 ( .A(n612), .B(n627), .CI(n610), .CO(n605), .S(n606) );
  CFA1X1 U502 ( .A(n631), .B(n629), .CI(n614), .CO(n607), .S(n608) );
  CFA1X1 U503 ( .A(n633), .B(n616), .CI(n618), .CO(n609), .S(n610) );
  CFA1X1 U504 ( .A(n635), .B(n620), .CI(n637), .CO(n611), .S(n612) );
  CFA1X1 U505 ( .A(n939), .B(n639), .CI(n622), .CO(n613), .S(n614) );
  CFA1X1 U507 ( .A(n901), .B(n1069), .CI(n985), .CO(n617), .S(n618) );
  CFA1X1 U508 ( .A(n859), .B(n1011), .CI(n871), .CO(n619), .S(n620) );
  CHA1X1 U509 ( .A(n808), .B(n885), .CO(n621), .S(n622) );
  CFA1X1 U511 ( .A(n632), .B(n645), .CI(n630), .CO(n625), .S(n626) );
  CFA1X1 U512 ( .A(n634), .B(n647), .CI(n649), .CO(n627), .S(n628) );
  CFA1X1 U513 ( .A(n640), .B(n636), .CI(n638), .CO(n629), .S(n630) );
  CFA1X1 U514 ( .A(n655), .B(n651), .CI(n653), .CO(n631), .S(n632) );
  CFA1X1 U515 ( .A(n940), .B(n657), .CI(n962), .CO(n633), .S(n634) );
  CFA1X1 U516 ( .A(n920), .B(n1040), .CI(n986), .CO(n635), .S(n636) );
  CFA1X1 U518 ( .A(n860), .B(n886), .CI(n872), .CO(n639), .S(n640) );
  CFA1X1 U519 ( .A(n646), .B(n644), .CI(n661), .CO(n641), .S(n642) );
  CFA1X1 U520 ( .A(n650), .B(n663), .CI(n648), .CO(n643), .S(n644) );
  CFA1X1 U521 ( .A(n652), .B(n665), .CI(n667), .CO(n645), .S(n646) );
  CFA1X1 U522 ( .A(n671), .B(n654), .CI(n656), .CO(n647), .S(n648) );
  CFA1X1 U523 ( .A(n658), .B(n669), .CI(n673), .CO(n649), .S(n650) );
  CFA1X1 U525 ( .A(n887), .B(n1041), .CI(n963), .CO(n653), .S(n654) );
  CFA1X1 U526 ( .A(n1071), .B(n873), .CI(n921), .CO(n655), .S(n656) );
  CHA1X1 U527 ( .A(n809), .B(n941), .CO(n657), .S(n658) );
  CFA1X1 U528 ( .A(n664), .B(n662), .CI(n677), .CO(n659), .S(n660) );
  CFA1X1 U529 ( .A(n668), .B(n679), .CI(n666), .CO(n661), .S(n662) );
  CFA1X1 U530 ( .A(n670), .B(n681), .CI(n683), .CO(n663), .S(n664) );
  CFA1X1 U532 ( .A(n964), .B(n687), .CI(n689), .CO(n667), .S(n668) );
  CFA1X1 U535 ( .A(n874), .B(n904), .CI(n888), .CO(n673), .S(n674) );
  CFA1X1 U538 ( .A(n688), .B(n697), .CI(n686), .CO(n679), .S(n680) );
  CFA1X1 U540 ( .A(n923), .B(n690), .CI(n943), .CO(n683), .S(n684) );
  CFA1X1 U541 ( .A(n905), .B(n1043), .CI(n1015), .CO(n685), .S(n686) );
  CFA1X1 U542 ( .A(n889), .B(n1073), .CI(n965), .CO(n687), .S(n688) );
  CFA1X1 U544 ( .A(n696), .B(n694), .CI(n707), .CO(n691), .S(n692) );
  CFA1X1 U545 ( .A(n711), .B(n709), .CI(n698), .CO(n693), .S(n694) );
  CFA1X1 U546 ( .A(n702), .B(n704), .CI(n700), .CO(n695), .S(n696) );
  CFA1X1 U547 ( .A(n717), .B(n715), .CI(n713), .CO(n697), .S(n698) );
  CFA1X1 U549 ( .A(n1074), .B(n1044), .CI(n944), .CO(n701), .S(n702) );
  CFA1X1 U550 ( .A(n890), .B(n906), .CI(n924), .CO(n703), .S(n704) );
  CFA1X1 U551 ( .A(n710), .B(n708), .CI(n721), .CO(n705), .S(n706) );
  CFA1X1 U552 ( .A(n725), .B(n723), .CI(n712), .CO(n707), .S(n708) );
  CFA1X1 U553 ( .A(n727), .B(n714), .CI(n716), .CO(n709), .S(n710) );
  CFA1X1 U554 ( .A(n945), .B(n729), .CI(n718), .CO(n711), .S(n712) );
  CFA1X1 U555 ( .A(n925), .B(n991), .CI(n967), .CO(n713), .S(n714) );
  CFA1X1 U556 ( .A(n1075), .B(n907), .CI(n1017), .CO(n715), .S(n716) );
  CFA1X1 U558 ( .A(n724), .B(n722), .CI(n733), .CO(n719), .S(n720) );
  CFA1X1 U559 ( .A(n728), .B(n735), .CI(n726), .CO(n721), .S(n722) );
  CFA1X1 U560 ( .A(n739), .B(n730), .CI(n737), .CO(n723), .S(n724) );
  CFA1X1 U561 ( .A(n992), .B(n741), .CI(n1630), .CO(n725), .S(n726) );
  CFA1X1 U562 ( .A(n968), .B(n1076), .CI(n1046), .CO(n727), .S(n728) );
  CFA1X1 U564 ( .A(n736), .B(n734), .CI(n745), .CO(n731), .S(n732) );
  CFA1X1 U565 ( .A(n740), .B(n747), .CI(n738), .CO(n733), .S(n734) );
  CFA1X1 U566 ( .A(n742), .B(n749), .CI(n751), .CO(n735), .S(n736) );
  CFA1X1 U567 ( .A(n993), .B(n947), .CI(n969), .CO(n737), .S(n738) );
  CFA1X1 U568 ( .A(n927), .B(n1047), .CI(n1019), .CO(n739), .S(n740) );
  CHA1X1 U569 ( .A(n812), .B(n1077), .CO(n741), .S(n742) );
  CFA1X1 U570 ( .A(n755), .B(n746), .CI(n748), .CO(n743), .S(n744) );
  CFA1X1 U571 ( .A(n752), .B(n757), .CI(n750), .CO(n745), .S(n746) );
  CFA1X1 U572 ( .A(n1020), .B(n759), .CI(n761), .CO(n747), .S(n748) );
  CFA1X1 U574 ( .A(n928), .B(n970), .CI(n948), .CO(n751), .S(n752) );
  CFA1X1 U575 ( .A(n758), .B(n756), .CI(n765), .CO(n753), .S(n754) );
  CFA1X1 U576 ( .A(n769), .B(n760), .CI(n767), .CO(n755), .S(n756) );
  CFA1X1 U577 ( .A(n971), .B(n762), .CI(n995), .CO(n757), .S(n758) );
  CFA1X1 U578 ( .A(n1049), .B(n949), .CI(n1021), .CO(n759), .S(n760) );
  CHA1X1 U579 ( .A(n813), .B(n1079), .CO(n761), .S(n762) );
  CFA1X1 U580 ( .A(n768), .B(n766), .CI(n773), .CO(n763), .S(n764) );
  CFA1X1 U581 ( .A(n777), .B(n770), .CI(n775), .CO(n765), .S(n766) );
  CFA1X1 U582 ( .A(n1022), .B(n1080), .CI(n1050), .CO(n767), .S(n768) );
  CFA1X1 U583 ( .A(n950), .B(n996), .CI(n972), .CO(n769), .S(n770) );
  CFA1X1 U584 ( .A(n781), .B(n774), .CI(n776), .CO(n771), .S(n772) );
  CFA1X1 U585 ( .A(n997), .B(n783), .CI(n778), .CO(n773), .S(n774) );
  CFA1X1 U586 ( .A(n973), .B(n1051), .CI(n1023), .CO(n775), .S(n776) );
  CHA1X1 U587 ( .A(n814), .B(n1081), .CO(n777), .S(n778) );
  CFA1X1 U588 ( .A(n787), .B(n782), .CI(n784), .CO(n779), .S(n780) );
  CFA1X1 U589 ( .A(n1052), .B(n789), .CI(n1082), .CO(n781), .S(n782) );
  CFA1X1 U591 ( .A(n790), .B(n788), .CI(n793), .CO(n785), .S(n786) );
  CFA1X1 U592 ( .A(n999), .B(n1053), .CI(n1025), .CO(n787), .S(n788) );
  CHA1X1 U593 ( .A(n815), .B(n1083), .CO(n789), .S(n790) );
  CFA1X1 U594 ( .A(n1084), .B(n794), .CI(n797), .CO(n791), .S(n792) );
  CFA1X1 U595 ( .A(n1000), .B(n1054), .CI(n1026), .CO(n793), .S(n794) );
  CFA1X1 U596 ( .A(n1027), .B(n798), .CI(n1055), .CO(n795), .S(n796) );
  CHA1X1 U597 ( .A(n816), .B(n1085), .CO(n797), .S(n798) );
  CFA1X1 U598 ( .A(n1028), .B(n1086), .CI(n1056), .CO(n799), .S(n800) );
  CHA1X1 U599 ( .A(n817), .B(n1057), .CO(n801), .S(n802) );
  COND2X1 U600 ( .A(n115), .B(n1435), .C(n114), .D(n1092), .Z(n803) );
  COND2X1 U601 ( .A(n1091), .B(n115), .C(n114), .D(n1090), .Z(n819) );
  COND2X1 U607 ( .A(n112), .B(n1094), .C(n110), .D(n1093), .Z(n821) );
  COND2X1 U608 ( .A(n112), .B(n1095), .C(n110), .D(n1094), .Z(n822) );
  COND2X1 U609 ( .A(n1096), .B(n112), .C(n110), .D(n1095), .Z(n823) );
  COND2X1 U620 ( .A(n107), .B(n1102), .C(n1101), .D(n105), .Z(n828) );
  COND2X1 U632 ( .A(n102), .B(n1107), .C(n1106), .D(n100), .Z(n832) );
  COND2X1 U635 ( .A(n102), .B(n1110), .C(n1109), .D(n100), .Z(n835) );
  COND2X1 U636 ( .A(n102), .B(n1111), .C(n1110), .D(n100), .Z(n836) );
  COND2X1 U637 ( .A(n1112), .B(n102), .C(n1111), .D(n100), .Z(n837) );
  COND2X1 U651 ( .A(n1565), .B(n1117), .C(n1116), .D(n95), .Z(n841) );
  COND2X1 U652 ( .A(n1565), .B(n1118), .C(n1117), .D(n1564), .Z(n842) );
  COND2X1 U655 ( .A(n97), .B(n1121), .C(n1120), .D(n95), .Z(n845) );
  COND2X1 U656 ( .A(n1565), .B(n1122), .C(n1121), .D(n1564), .Z(n846) );
  COND2X1 U657 ( .A(n1565), .B(n1123), .C(n1122), .D(n1564), .Z(n847) );
  COND2X1 U670 ( .A(n1572), .B(n1871), .C(n1137), .D(n1650), .Z(n808) );
  COND2X1 U677 ( .A(n1572), .B(n1132), .C(n1131), .D(n1650), .Z(n855) );
  COND2X1 U680 ( .A(n1572), .B(n1135), .C(n1134), .D(n1651), .Z(n858) );
  COND2X1 U681 ( .A(n1572), .B(n1136), .C(n1135), .D(n1651), .Z(n859) );
  COND2X1 U696 ( .A(n84), .B(n1866), .C(n1152), .D(n1781), .Z(n809) );
  COND2X1 U697 ( .A(n84), .B(n1139), .C(n1138), .D(n1781), .Z(n861) );
  COND2X1 U698 ( .A(n84), .B(n1140), .C(n1139), .D(n1781), .Z(n862) );
  COND2X1 U699 ( .A(n84), .B(n1141), .C(n1140), .D(n1781), .Z(n863) );
  COND2X1 U701 ( .A(n84), .B(n1143), .C(n1142), .D(n1781), .Z(n865) );
  COND2X1 U702 ( .A(n84), .B(n1144), .C(n1143), .D(n1781), .Z(n866) );
  COND2X1 U703 ( .A(n84), .B(n1145), .C(n1144), .D(n1781), .Z(n867) );
  COND2X1 U707 ( .A(n84), .B(n1149), .C(n1148), .D(n1781), .Z(n871) );
  COND2X1 U708 ( .A(n84), .B(n1150), .C(n1149), .D(n1781), .Z(n872) );
  COND2X1 U709 ( .A(n84), .B(n1151), .C(n1150), .D(n1781), .Z(n873) );
  COND2X1 U728 ( .A(n77), .B(n1155), .C(n1154), .D(n1638), .Z(n876) );
  COND2X1 U729 ( .A(n77), .B(n1156), .C(n1155), .D(n1638), .Z(n877) );
  COND2X1 U730 ( .A(n77), .B(n1157), .C(n1156), .D(n1638), .Z(n878) );
  COND2X1 U731 ( .A(n77), .B(n1158), .C(n1157), .D(n1638), .Z(n879) );
  COND2X1 U732 ( .A(n77), .B(n1159), .C(n1158), .D(n1639), .Z(n880) );
  COND2X1 U733 ( .A(n77), .B(n1160), .C(n1159), .D(n1638), .Z(n881) );
  COND2X1 U734 ( .A(n77), .B(n1161), .C(n1160), .D(n1639), .Z(n882) );
  COND2X1 U735 ( .A(n77), .B(n1162), .C(n1161), .D(n1638), .Z(n883) );
  COND2X1 U737 ( .A(n77), .B(n1164), .C(n1163), .D(n1639), .Z(n885) );
  COND2X1 U738 ( .A(n77), .B(n1165), .C(n1164), .D(n1639), .Z(n886) );
  COND2X1 U739 ( .A(n77), .B(n1166), .C(n1165), .D(n1639), .Z(n887) );
  COND2X1 U741 ( .A(n77), .B(n1168), .C(n1167), .D(n1639), .Z(n889) );
  COND2X1 U764 ( .A(n69), .B(n1174), .C(n1173), .D(n1776), .Z(n894) );
  COND2X1 U765 ( .A(n69), .B(n1175), .C(n1174), .D(n1777), .Z(n895) );
  COND2X1 U766 ( .A(n69), .B(n1176), .C(n1175), .D(n1777), .Z(n896) );
  COND2X1 U767 ( .A(n69), .B(n1177), .C(n1176), .D(n1776), .Z(n897) );
  COND2X1 U768 ( .A(n69), .B(n1178), .C(n1177), .D(n1776), .Z(n898) );
  COND2X1 U771 ( .A(n69), .B(n1181), .C(n1180), .D(n1777), .Z(n901) );
  COND2X1 U775 ( .A(n69), .B(n1185), .C(n1184), .D(n1777), .Z(n905) );
  COND2X1 U803 ( .A(n61), .B(n1194), .C(n1193), .D(n58), .Z(n913) );
  COND2X1 U804 ( .A(n1195), .B(n61), .C(n1194), .D(n58), .Z(n914) );
  COND2X1 U805 ( .A(n61), .B(n1196), .C(n1195), .D(n58), .Z(n915) );
  COND2X1 U811 ( .A(n61), .B(n1202), .C(n1201), .D(n58), .Z(n921) );
  COND2X1 U812 ( .A(n61), .B(n1203), .C(n1202), .D(n58), .Z(n922) );
  COND2X1 U814 ( .A(n61), .B(n1205), .C(n1204), .D(n58), .Z(n924) );
  COND2X1 U815 ( .A(n61), .B(n1206), .C(n1205), .D(n58), .Z(n925) );
  COND2X1 U816 ( .A(n61), .B(n1207), .C(n1206), .D(n58), .Z(n926) );
  COND2X1 U847 ( .A(n53), .B(n1217), .C(n1216), .D(n50), .Z(n935) );
  COND2X1 U856 ( .A(n1559), .B(n1226), .C(n1225), .D(n50), .Z(n944) );
  COND2X1 U886 ( .A(n1653), .B(n1845), .C(n1257), .D(n1576), .Z(n814) );
  COND2X1 U890 ( .A(n1654), .B(n1237), .C(n1236), .D(n1575), .Z(n954) );
  COND2X1 U892 ( .A(n1654), .B(n1239), .C(n1238), .D(n1575), .Z(n956) );
  COND2X1 U893 ( .A(n1654), .B(n1240), .C(n1239), .D(n1575), .Z(n957) );
  COND2X1 U894 ( .A(n1653), .B(n1241), .C(n1240), .D(n1575), .Z(n958) );
  COND2X1 U897 ( .A(n1653), .B(n1244), .C(n1243), .D(n1575), .Z(n961) );
  COND2X1 U899 ( .A(n1653), .B(n1246), .C(n1245), .D(n1575), .Z(n963) );
  COND2X1 U901 ( .A(n1653), .B(n1248), .C(n1247), .D(n1576), .Z(n965) );
  COND2X1 U904 ( .A(n1654), .B(n1251), .C(n1250), .D(n1576), .Z(n968) );
  COND2X1 U905 ( .A(n1654), .B(n1252), .C(n1251), .D(n1575), .Z(n969) );
  COND2X1 U906 ( .A(n1654), .B(n1253), .C(n1252), .D(n1576), .Z(n970) );
  COND2X1 U908 ( .A(n1653), .B(n1255), .C(n1254), .D(n1575), .Z(n972) );
  COND2X1 U909 ( .A(n1654), .B(n1256), .C(n1255), .D(n1575), .Z(n973) );
  CND2IX1 U935 ( .B(n1876), .A(n1839), .Z(n1257) );
  COND2X1 U941 ( .A(n1571), .B(n1263), .C(n1262), .D(n1796), .Z(n979) );
  COND2X1 U942 ( .A(n36), .B(n1264), .C(n1263), .D(n1796), .Z(n980) );
  COND2X1 U943 ( .A(n36), .B(n1265), .C(n1264), .D(n1796), .Z(n981) );
  COND2X1 U944 ( .A(n1570), .B(n1266), .C(n1265), .D(n1796), .Z(n982) );
  COND2X1 U946 ( .A(n1570), .B(n1268), .C(n1267), .D(n1796), .Z(n984) );
  COND2X1 U947 ( .A(n1571), .B(n1269), .C(n1268), .D(n1796), .Z(n985) );
  COND2X1 U948 ( .A(n1571), .B(n1270), .C(n1269), .D(n1796), .Z(n986) );
  COND2X1 U952 ( .A(n1571), .B(n1274), .C(n1273), .D(n1796), .Z(n990) );
  COND2X1 U953 ( .A(n1570), .B(n1275), .C(n1274), .D(n1796), .Z(n991) );
  COND2X1 U958 ( .A(n1570), .B(n1280), .C(n1279), .D(n1796), .Z(n996) );
  COND2X1 U992 ( .A(n1619), .B(n1287), .C(n1286), .D(n24), .Z(n1002) );
  COND2X1 U993 ( .A(n1619), .B(n1288), .C(n1287), .D(n24), .Z(n1003) );
  COND2X1 U995 ( .A(n1619), .B(n1290), .C(n1289), .D(n24), .Z(n1005) );
  COND2X1 U996 ( .A(n27), .B(n1291), .C(n1290), .D(n24), .Z(n1006) );
  COND2X1 U997 ( .A(n1620), .B(n1292), .C(n1291), .D(n24), .Z(n1007) );
  COND2X1 U1000 ( .A(n1619), .B(n1295), .C(n1294), .D(n24), .Z(n1010) );
  COND2X1 U1001 ( .A(n1620), .B(n1296), .C(n1295), .D(n24), .Z(n1011) );
  COND2X1 U1002 ( .A(n1619), .B(n1297), .C(n1296), .D(n24), .Z(n1012) );
  COND2X1 U1005 ( .A(n1619), .B(n1300), .C(n1299), .D(n24), .Z(n1015) );
  COND2X1 U1006 ( .A(n1619), .B(n1301), .C(n1300), .D(n24), .Z(n1016) );
  COND2X1 U1007 ( .A(n27), .B(n1302), .C(n1301), .D(n24), .Z(n1017) );
  COND2X1 U1009 ( .A(n1620), .B(n1304), .C(n1303), .D(n24), .Z(n1019) );
  COND2X1 U1011 ( .A(n1620), .B(n1306), .C(n1305), .D(n24), .Z(n1021) );
  COND2X1 U1012 ( .A(n1620), .B(n1307), .C(n1306), .D(n24), .Z(n1022) );
  COND2X1 U1013 ( .A(n1619), .B(n1308), .C(n1307), .D(n24), .Z(n1023) );
  COND2X1 U1016 ( .A(n1620), .B(n1311), .C(n1310), .D(n24), .Z(n1026) );
  CND2IX1 U1047 ( .B(n1876), .A(n1588), .Z(n1313) );
  COND2X1 U1051 ( .A(n18), .B(n1317), .C(n1316), .D(n1574), .Z(n1031) );
  COND2X1 U1052 ( .A(n18), .B(n1318), .C(n1317), .D(n1574), .Z(n1032) );
  COND2X1 U1053 ( .A(n18), .B(n1319), .C(n1318), .D(n1574), .Z(n1033) );
  COND2X1 U1054 ( .A(n18), .B(n1320), .C(n1319), .D(n1573), .Z(n1034) );
  COND2X1 U1055 ( .A(n18), .B(n1321), .C(n1320), .D(n1574), .Z(n1035) );
  COND2X1 U1056 ( .A(n18), .B(n1322), .C(n1321), .D(n1573), .Z(n1036) );
  COND2X1 U1061 ( .A(n18), .B(n1327), .C(n1326), .D(n1574), .Z(n1041) );
  COND2X1 U1062 ( .A(n18), .B(n1328), .C(n1327), .D(n1574), .Z(n1042) );
  COND2X1 U1064 ( .A(n18), .B(n1330), .C(n1329), .D(n1574), .Z(n1044) );
  COND2X1 U1065 ( .A(n18), .B(n1331), .C(n1330), .D(n1573), .Z(n1045) );
  COND2X1 U1066 ( .A(n18), .B(n1332), .C(n1331), .D(n1573), .Z(n1046) );
  COND2X1 U1067 ( .A(n18), .B(n1333), .C(n1332), .D(n1574), .Z(n1047) );
  COND2X1 U1068 ( .A(n18), .B(n1334), .C(n1333), .D(n1573), .Z(n1048) );
  COND2X1 U1069 ( .A(n18), .B(n1335), .C(n1334), .D(n1574), .Z(n1049) );
  COND2X1 U1071 ( .A(n18), .B(n1337), .C(n1336), .D(n1573), .Z(n1051) );
  COND2X1 U1074 ( .A(n18), .B(n1340), .C(n1339), .D(n1573), .Z(n1054) );
  CEOX2 U1261 ( .A(a[4]), .B(n1829), .Z(n1423) );
  CFD1QX1 clk_r_REG312_S1 ( .D(n1705), .CP(n1774), .Q(n1773) );
  CFD1QX1 clk_r_REG319_S1 ( .D(n355), .CP(n1774), .Q(n1771) );
  CFD1QX1 clk_r_REG311_S1 ( .D(n256), .CP(n1774), .Q(n1770) );
  CFD1QX1 clk_r_REG310_S1 ( .D(n258), .CP(n1774), .Q(n1769) );
  CFD1QX1 clk_r_REG318_S1 ( .D(n281), .CP(n1774), .Q(n1764) );
  CFD1QX1 clk_r_REG289_S1 ( .D(n284), .CP(n1774), .Q(n1763) );
  CFD1QX1 clk_r_REG286_S1 ( .D(n290), .CP(n1774), .Q(n1760) );
  CFD1QX1 clk_r_REG285_S1 ( .D(n140), .CP(n1774), .Q(n1759) );
  CFD1QX1 clk_r_REG328_S1 ( .D(n1799), .CP(n1774), .Q(n1758) );
  CFD1QX1 clk_r_REG299_S1 ( .D(n441), .CP(n1774), .Q(n1745) );
  CFD1QX1 clk_r_REG298_S1 ( .D(n444), .CP(n1774), .Q(n1743) );
  CFD1QX1 clk_r_REG296_S1 ( .D(n467), .CP(n1774), .Q(n1742) );
  CFD1QX1 clk_r_REG297_S1 ( .D(n468), .CP(n1774), .Q(n1741) );
  CFD1QX1 clk_r_REG335_S1 ( .D(n470), .CP(n1774), .Q(n1740) );
  CFD1QX1 clk_r_REG333_S1 ( .D(n493), .CP(n1774), .Q(n1739) );
  CFD1QX1 clk_r_REG334_S1 ( .D(n494), .CP(n1774), .Q(n1738) );
  CFD1QX1 clk_r_REG343_S1 ( .D(n496), .CP(n1774), .Q(n1737) );
  CFD1QX1 clk_r_REG336_S1 ( .D(n517), .CP(n1774), .Q(n1736) );
  CFD1QX1 clk_r_REG337_S1 ( .D(n518), .CP(n1774), .Q(n1735) );
  CFD1QX1 clk_r_REG332_S1 ( .D(n520), .CP(n1774), .Q(n1734) );
  CFD1QX1 clk_r_REG329_S1 ( .D(n541), .CP(n1774), .Q(n1733) );
  CFD1QX1 clk_r_REG330_S1 ( .D(n542), .CP(n1774), .Q(n1732) );
  CFD1QX1 clk_r_REG326_S1 ( .D(n563), .CP(n1774), .Q(n1730) );
  CFD1QX1 clk_r_REG327_S1 ( .D(n564), .CP(n1774), .Q(net171532) );
  CFD1QX1 clk_r_REG324_S1 ( .D(n606), .CP(n1774), .Q(net171538) );
  CFD1QX1 clk_r_REG316_S1 ( .D(n641), .CP(n1774), .Q(n1727) );
  CFD1QX1 clk_r_REG317_S1 ( .D(n642), .CP(n1774), .Q(n1726) );
  CFD1QX1 clk_r_REG314_S1 ( .D(n659), .CP(n1774), .Q(n1724) );
  CFD1QX1 clk_r_REG315_S1 ( .D(n660), .CP(n1774), .Q(n1723) );
  CFD1QX1 clk_r_REG313_S1 ( .D(n675), .CP(n1774), .Q(n1722) );
  CFD1QXL clk_r_REG302_S1 ( .D(n385), .CP(n1774), .Q(n1752) );
  CFD1QXL clk_r_REG293_S1 ( .D(n369), .CP(n1774), .Q(n1755) );
  CFD1QXL clk_r_REG294_S1 ( .D(n413), .CP(n1774), .Q(n1748) );
  CFD1QXL clk_r_REG292_S1 ( .D(n388), .CP(n1774), .Q(n1749) );
  CFD1QX4 clk_r_REG322_S1 ( .D(n626), .CP(n1774), .Q(n1729) );
  CFD1QX2 clk_r_REG331_S1 ( .D(n628), .CP(n1774), .Q(n1728) );
  CFD1QX4 clk_r_REG325_S1 ( .D(n588), .CP(n1774), .Q(net171536) );
  CFD1QX2 clk_r_REG287_S1 ( .D(n285), .CP(n1774), .Q(n1757) );
  CFD1QX2 clk_r_REG339_S1 ( .D(n585), .CP(n1774), .Q(net171534) );
  CFD1QX2 clk_r_REG321_S1 ( .D(n625), .CP(n1774), .Q(net171540) );
  CFD1QX2 clk_r_REG308_S1 ( .D(n1706), .CP(n1774), .Q(n1772) );
  CFD1QX2 clk_r_REG283_S1 ( .D(n292), .CP(n1774), .Q(n1754) );
  CFD1QX2 clk_r_REG288_S1 ( .D(n289), .CP(n1774), .Q(n1761) );
  CFD1QX4 clk_r_REG320_S1 ( .D(n643), .CP(n1774), .Q(n1725) );
  CFD1QX2 clk_r_REG307_S1 ( .D(n271), .CP(n1774), .Q(n1767) );
  CFD1QX2 clk_r_REG306_S1 ( .D(n273), .CP(n1774), .Q(n1766) );
  CFD1QX2 clk_r_REG304_S1 ( .D(n136), .CP(n1774), .Q(n1765) );
  CFD1QX2 clk_r_REG309_S1 ( .D(n259), .CP(n1774), .Q(n1768) );
  CFD1QX2 clk_r_REG284_S1 ( .D(n299), .CP(n1774), .Q(n1756) );
  CFD1QX2 clk_r_REG290_S1 ( .D(n138), .CP(n1774), .Q(n1762) );
  CFA1X1 U479 ( .A(net171533), .B(net171532), .CI(net171534), .CO(n561), .S(
        n562) );
  CANR1X1 U123 ( .A(n182), .B(n169), .C(n170), .Z(n168) );
  COND1X1 U125 ( .A(n179), .B(n171), .C(n172), .Z(n170) );
  CNR2X2 U197 ( .A(net179596), .B(n603), .Z(n222) );
  CFA1X1 U500 ( .A(net171539), .B(net171538), .CI(net171540), .CO(n603), .S(
        n604) );
  CFA1X1 U490 ( .A(net171536), .B(net171535), .CI(net171537), .CO(n583), .S(
        n584) );
  CFD1QXL clk_r_REG301_S1 ( .D(n416), .CP(n1774), .Q(n1746) );
  CFD1QXL clk_r_REG291_S1 ( .D(n387), .CP(n1774), .Q(n1750) );
  CFD1QXL clk_r_REG342_S1 ( .D(n544), .CP(n1774), .Q(n1731) );
  CFD1QX2 clk_r_REG305_S1 ( .D(n274), .CP(n1774), .Q(n1753) );
  CFD1QX2 clk_r_REG338_S1 ( .D(n608), .CP(n1774), .Q(net171539) );
  CFD1QX2 clk_r_REG323_S1 ( .D(n605), .CP(n1774), .Q(net171537) );
  CFD1QX4 clk_r_REG341_S1 ( .D(n566), .CP(n1774), .Q(net171533) );
  CFD1QX2 clk_r_REG295_S1 ( .D(n414), .CP(n1774), .Q(n1747) );
  CFD1QX2 clk_r_REG303_S1 ( .D(n386), .CP(n1774), .Q(n1751) );
  CFD1QX2 clk_r_REG300_S1 ( .D(n442), .CP(n1774), .Q(n1744) );
  CFD1QX2 clk_r_REG340_S1 ( .D(n586), .CP(n1774), .Q(net171535) );
  CNR2X2 U1271 ( .A(n6), .B(n1349), .Z(n1063) );
  CNR2X2 U1272 ( .A(n6), .B(n1351), .Z(n1065) );
  CNR2X2 U1273 ( .A(n6), .B(n1361), .Z(n1075) );
  CNR2X2 U1274 ( .A(n6), .B(n1360), .Z(n1074) );
  CNR2X2 U1275 ( .A(n6), .B(n1358), .Z(n1072) );
  CNR2X2 U1276 ( .A(n6), .B(n1357), .Z(n1071) );
  CNR2X2 U1277 ( .A(n6), .B(n1348), .Z(n1062) );
  CNR2X2 U1278 ( .A(n6), .B(n1363), .Z(n1077) );
  CNR2X2 U1279 ( .A(n6), .B(n1350), .Z(n1064) );
  CNR2X2 U1280 ( .A(n6), .B(n1374), .Z(n1088) );
  CNR2X2 U1281 ( .A(n6), .B(n1364), .Z(n1078) );
  CNR2X2 U1282 ( .A(n6), .B(n1354), .Z(n1068) );
  CNR2X2 U1283 ( .A(n6), .B(n1347), .Z(n1061) );
  CNR2X2 U1284 ( .A(n6), .B(n1365), .Z(n1079) );
  CNR2X2 U1285 ( .A(n6), .B(n1359), .Z(n1073) );
  CNR2X2 U1286 ( .A(n6), .B(n1355), .Z(n1069) );
  CNR2X2 U1287 ( .A(n6), .B(n1352), .Z(n1066) );
  CNR2X2 U1288 ( .A(n6), .B(n1369), .Z(n1083) );
  CNR2X2 U1289 ( .A(n6), .B(n1371), .Z(n1085) );
  CNR2X2 U1290 ( .A(n6), .B(n1362), .Z(n1076) );
  CNR2X2 U1291 ( .A(n6), .B(n1367), .Z(n1081) );
  CNR2X2 U1292 ( .A(n6), .B(n1372), .Z(n1086) );
  CNR2X2 U1293 ( .A(n6), .B(n1353), .Z(n1067) );
  CNR2X2 U1294 ( .A(n6), .B(n1356), .Z(n1070) );
  CNR2X2 U1295 ( .A(n6), .B(n1368), .Z(n1082) );
  CNR2X2 U1296 ( .A(n6), .B(n1346), .Z(n1060) );
  CNR2X2 U1297 ( .A(n6), .B(n1366), .Z(n1080) );
  CNR2X2 U1298 ( .A(n6), .B(n1370), .Z(n1084) );
  CNR2X2 U1299 ( .A(n6), .B(n1373), .Z(n1087) );
  CNR2X2 U1300 ( .A(n6), .B(n1345), .Z(n1059) );
  CNR2X2 U1301 ( .A(n6), .B(n1375), .Z(n1089) );
  CIVX2 U1302 ( .A(a[2]), .Z(n1590) );
  CIVX2 U1303 ( .A(a[2]), .Z(n1573) );
  CIVX2 U1304 ( .A(a[2]), .Z(n1574) );
  CIVX2 U1305 ( .A(n1393), .Z(n1360) );
  CIVX2 U1306 ( .A(n1817), .Z(n1362) );
  CIVX2 U1307 ( .A(n1818), .Z(n1361) );
  CIVX2 U1308 ( .A(n1815), .Z(n1364) );
  CIVX2 U1309 ( .A(n1392), .Z(n1359) );
  CIVX2 U1310 ( .A(n1816), .Z(n1363) );
  CIVX2 U1311 ( .A(n1089), .Z(n335) );
  CIVX2 U1312 ( .A(n335), .Z(product[1]) );
  CIVX2 U1313 ( .A(n148), .Z(product[2]) );
  CIVX2 U1314 ( .A(n331), .Z(n329) );
  CIVX2 U1315 ( .A(n1388), .Z(n1355) );
  CIVX2 U1316 ( .A(n1386), .Z(n1353) );
  CIVX2 U1317 ( .A(n1390), .Z(n1357) );
  CIVX2 U1318 ( .A(n1389), .Z(n1356) );
  CIVX2 U1319 ( .A(b[25]), .Z(n1351) );
  CIVX2 U1320 ( .A(b[24]), .Z(n1352) );
  CIVX2 U1321 ( .A(b[28]), .Z(n1348) );
  CIVX2 U1322 ( .A(b[30]), .Z(n1346) );
  CIVX2 U1323 ( .A(n1811), .Z(n1369) );
  CIVX2 U1324 ( .A(b[29]), .Z(n1347) );
  CIVX2 U1325 ( .A(b[26]), .Z(n1350) );
  CIVX2 U1326 ( .A(n1387), .Z(n1354) );
  CIVX2 U1327 ( .A(b[27]), .Z(n1349) );
  CIVX2 U1328 ( .A(b[31]), .Z(n1345) );
  CIVX2 U1329 ( .A(n1807), .Z(n1373) );
  CIVX2 U1330 ( .A(n1813), .Z(n1366) );
  CIVX2 U1331 ( .A(n1810), .Z(n1370) );
  CIVX2 U1332 ( .A(n1806), .Z(n1374) );
  CIVX2 U1333 ( .A(n1805), .Z(n1375) );
  CIVX2 U1334 ( .A(n1814), .Z(n1365) );
  CIVX2 U1335 ( .A(n1401), .Z(n1368) );
  CIVX2 U1336 ( .A(n1391), .Z(n1358) );
  CIVX2 U1337 ( .A(n1812), .Z(n1367) );
  CIVX2 U1338 ( .A(n1808), .Z(n1372) );
  CIVX2 U1339 ( .A(n1809), .Z(n1371) );
  COAN1X1 U1340 ( .A(n233), .B(n245), .C(n234), .Z(n1549) );
  CIVX1 U1341 ( .A(n1551), .Z(net179577) );
  COND1X1 U1342 ( .A(n198), .B(n1548), .C(n199), .Z(n1547) );
  CANR1X1 U1343 ( .A(n228), .B(n346), .C(n1581), .Z(n1548) );
  COND1X1 U1344 ( .A(n198), .B(n215), .C(n199), .Z(n197) );
  CANR1X1 U1345 ( .A(n228), .B(n346), .C(n1581), .Z(n215) );
  CIVXL U1346 ( .A(n222), .Z(n1550) );
  CAOR1X1 U1347 ( .A(n228), .B(n1550), .C(net179873), .Z(n1551) );
  CND2X2 U1348 ( .A(n348), .B(n349), .Z(n233) );
  CND2X1 U1349 ( .A(n1673), .B(net180181), .Z(n1554) );
  CND2X2 U1350 ( .A(n1552), .B(n1553), .Z(n1555) );
  CND2X2 U1351 ( .A(n1554), .B(n1555), .Z(product[22]) );
  CIVX2 U1352 ( .A(n1673), .Z(n1552) );
  CIVX2 U1353 ( .A(net180181), .Z(n1553) );
  CANR1X2 U1354 ( .A(net178506), .B(n166), .C(n163), .Z(n1625) );
  CENX2 U1355 ( .A(n1624), .B(n1625), .Z(product[30]) );
  CIVX1 U1356 ( .A(n298), .Z(n296) );
  CIVX1 U1357 ( .A(n50), .Z(n1556) );
  CIVX1 U1358 ( .A(n1556), .Z(n1557) );
  CND2IX2 U1359 ( .B(n1720), .A(n50), .Z(n1558) );
  CND2IX2 U1360 ( .B(n1720), .A(n50), .Z(n1559) );
  CND2IX1 U1361 ( .B(n1720), .A(n50), .Z(n53) );
  CNIVX1 U1362 ( .A(n50), .Z(n1560) );
  CENX1 U1363 ( .A(n1561), .B(n264), .Z(product[16]) );
  CAN2X2 U1364 ( .A(n352), .B(n1768), .Z(n1561) );
  CIVX1 U1365 ( .A(n934), .Z(n1562) );
  CIVX2 U1366 ( .A(n1562), .Z(n1563) );
  CIVX2 U1367 ( .A(n265), .Z(n264) );
  CEOX1 U1368 ( .A(n1631), .B(n454), .Z(n446) );
  CND2XL U1369 ( .A(n452), .B(n454), .Z(n1636) );
  COND2XL U1370 ( .A(n1103), .B(n107), .C(n105), .D(n1102), .Z(n829) );
  CNIVX4 U1371 ( .A(n95), .Z(n1564) );
  CND2X2 U1372 ( .A(n1414), .B(n95), .Z(n1565) );
  CND2X1 U1373 ( .A(n1414), .B(n95), .Z(n97) );
  COND2X1 U1374 ( .A(n84), .B(n1146), .C(n1145), .D(n1781), .Z(n868) );
  COND2XL U1375 ( .A(n84), .B(n1147), .C(n1146), .D(n1781), .Z(n869) );
  COND2XL U1376 ( .A(n84), .B(n1142), .C(n1141), .D(n1781), .Z(n864) );
  CIVXL U1377 ( .A(n55), .Z(n1566) );
  COND2X1 U1378 ( .A(n1654), .B(n1243), .C(n1242), .D(n1576), .Z(n960) );
  CENX2 U1379 ( .A(a[10]), .B(n1848), .Z(n1720) );
  CIVX2 U1380 ( .A(n1679), .Z(n1567) );
  CIVX1 U1381 ( .A(n1679), .Z(n1678) );
  COND2XL U1382 ( .A(n1565), .B(n1784), .C(n95), .D(n1124), .Z(n807) );
  CIVX1 U1383 ( .A(n1770), .Z(n254) );
  CIVX4 U1384 ( .A(n1850), .Z(n1848) );
  CIVXL U1385 ( .A(n1824), .Z(n1568) );
  CENX1 U1386 ( .A(a[12]), .B(n1566), .Z(n1419) );
  CENX1 U1387 ( .A(n1569), .B(n432), .Z(n422) );
  CENX1 U1388 ( .A(n430), .B(n434), .Z(n1569) );
  CNIVX4 U1389 ( .A(n1396), .Z(n1816) );
  CIVX4 U1390 ( .A(n1621), .Z(n1869) );
  CIVX4 U1391 ( .A(n1868), .Z(n1621) );
  CIVX1 U1392 ( .A(n1704), .Z(n1781) );
  COND2XL U1393 ( .A(n77), .B(n1163), .C(n1162), .D(n1638), .Z(n884) );
  COND2XL U1394 ( .A(n77), .B(n1154), .C(n1153), .D(n1639), .Z(n875) );
  CIVX3 U1395 ( .A(n1847), .Z(n1844) );
  CND2X2 U1396 ( .A(n1421), .B(n1804), .Z(n1653) );
  CENXL U1397 ( .A(n1842), .B(n1814), .Z(n1245) );
  CEOX2 U1398 ( .A(n1832), .B(a[6]), .Z(n33) );
  CND2X2 U1399 ( .A(n1422), .B(n1803), .Z(n1570) );
  CND2X2 U1400 ( .A(n1422), .B(n1803), .Z(n1571) );
  CND2X1 U1401 ( .A(n1422), .B(n1803), .Z(n36) );
  CANR1X2 U1402 ( .A(n318), .B(n1712), .C(n315), .Z(n313) );
  CNIVX4 U1403 ( .A(n33), .Z(n1803) );
  CENX1 U1404 ( .A(a[20]), .B(n1872), .Z(n1699) );
  CND2X2 U1405 ( .A(n1699), .B(n89), .Z(n1572) );
  CND2XL U1406 ( .A(n1699), .B(n89), .Z(n91) );
  CNIVX4 U1407 ( .A(n42), .Z(n1575) );
  CNIVX4 U1408 ( .A(n42), .Z(n1576) );
  CNIVX2 U1409 ( .A(n42), .Z(n1804) );
  CENXL U1410 ( .A(n1819), .B(b[29]), .Z(n1314) );
  CENXL U1411 ( .A(n1822), .B(n1814), .Z(n1332) );
  CNIVX1 U1412 ( .A(n833), .Z(n1577) );
  CENXL U1413 ( .A(n142), .B(n310), .Z(product[8]) );
  CENXL U1414 ( .A(n1822), .B(n1388), .Z(n1322) );
  CFA1XL U1415 ( .A(n917), .B(n1067), .CI(n1037), .CO(n575), .S(n576) );
  CND2X1 U1416 ( .A(net178515), .B(net178516), .Z(n1578) );
  CIVX1 U1417 ( .A(n305), .Z(n304) );
  CENX2 U1418 ( .A(n1579), .B(n1701), .Z(product[14]) );
  CIVX20 U1419 ( .A(n1765), .Z(n1579) );
  CHA1X1 U1420 ( .A(n810), .B(n989), .CO(n689), .S(n690) );
  CENXL U1421 ( .A(n1836), .B(n1814), .Z(n1272) );
  CND3X1 U1422 ( .A(n1666), .B(n1667), .C(n1668), .Z(n459) );
  CND2X1 U1423 ( .A(n357), .B(n1760), .Z(n1580) );
  CIVX3 U1424 ( .A(n1761), .Z(n357) );
  CENX1 U1425 ( .A(n1860), .B(n1816), .Z(n1155) );
  CIVX2 U1426 ( .A(net179871), .Z(n1581) );
  CIVXL U1427 ( .A(net179871), .Z(net179873) );
  COND1X1 U1428 ( .A(n167), .B(net181713), .C(n168), .Z(n166) );
  CAN2X1 U1429 ( .A(net178510), .B(n160), .Z(n1624) );
  CND2XL U1430 ( .A(n485), .B(n487), .Z(n1634) );
  CIVX3 U1431 ( .A(n1832), .Z(n1829) );
  CNR2X1 U1432 ( .A(n440), .B(n465), .Z(n171) );
  CND2X1 U1433 ( .A(n466), .B(n491), .Z(n179) );
  CIVX2 U1434 ( .A(n1867), .Z(n1865) );
  CIVX3 U1435 ( .A(n1866), .Z(n1862) );
  CENX1 U1436 ( .A(n1873), .B(n1808), .Z(n1108) );
  CND2X1 U1437 ( .A(n492), .B(n515), .Z(n188) );
  CND2X1 U1438 ( .A(n1726), .B(n1724), .Z(n243) );
  CENX1 U1439 ( .A(n1596), .B(n674), .Z(n666) );
  CENX1 U1440 ( .A(n685), .B(n672), .Z(n1596) );
  CND2XL U1441 ( .A(n489), .B(n485), .Z(n1632) );
  CIVX2 U1442 ( .A(n1587), .Z(n1831) );
  CIVDX2 U1443 ( .A(n55), .Z0(n1582), .Z1(n1583) );
  CIVDX1 U1444 ( .A(n30), .Z0(n1584), .Z1(n1585) );
  CNR2X1 U1445 ( .A(n150), .B(n1718), .Z(n1586) );
  CIVDX1 U1446 ( .A(n21), .Z0(n1587), .Z1(n1588) );
  CIVX2 U1447 ( .A(n1847), .Z(n1843) );
  CNIVX1 U1448 ( .A(n1038), .Z(n1589) );
  CIVX2 U1449 ( .A(net180264), .Z(net180393) );
  CAN2XL U1450 ( .A(n216), .B(net180512), .Z(n1591) );
  CAN2XL U1451 ( .A(net178510), .B(net178506), .Z(n1592) );
  CIVXL U1452 ( .A(n1437), .Z(n1593) );
  COR2XL U1453 ( .A(n772), .B(n779), .Z(n1594) );
  CIVX4 U1454 ( .A(n1595), .Z(n1849) );
  CND2X2 U1455 ( .A(n1707), .B(n303), .Z(n141) );
  COND2XL U1456 ( .A(n1565), .B(n1115), .C(n1114), .D(n1564), .Z(n839) );
  CND2IXL U1457 ( .B(n1876), .A(n93), .Z(n1124) );
  CENXL U1458 ( .A(n93), .B(n1806), .Z(n1121) );
  COND2XL U1459 ( .A(n97), .B(n1119), .C(n1118), .D(n95), .Z(n843) );
  CIVX1 U1460 ( .A(n48), .Z(n1595) );
  CIVX2 U1461 ( .A(n48), .Z(n1850) );
  CENX1 U1462 ( .A(n1869), .B(n1807), .Z(n1133) );
  COND2XL U1463 ( .A(n91), .B(n1133), .C(n1132), .D(n1650), .Z(n856) );
  CIVX2 U1464 ( .A(n1856), .Z(n1855) );
  CND2IX1 U1465 ( .B(n129), .A(n1549), .Z(n1656) );
  COND2X1 U1466 ( .A(n61), .B(n1788), .C(n1209), .D(n58), .Z(n812) );
  CIVXL U1467 ( .A(n113), .Z(n1435) );
  CIVX1 U1468 ( .A(n1861), .Z(n1858) );
  CIVX1 U1469 ( .A(n1861), .Z(n1860) );
  CIVX1 U1470 ( .A(n79), .Z(n1866) );
  CIVX3 U1471 ( .A(n1584), .Z(n1837) );
  CIVX2 U1472 ( .A(n21), .Z(n1832) );
  CENXL U1473 ( .A(n1865), .B(n1816), .Z(n1138) );
  CENXL U1474 ( .A(n1842), .B(n1816), .Z(n1243) );
  CENXL U1475 ( .A(n1854), .B(n1816), .Z(n1174) );
  COND2X1 U1476 ( .A(n1565), .B(n1116), .C(n1115), .D(n95), .Z(n840) );
  CND2X1 U1477 ( .A(n720), .B(n731), .Z(n276) );
  COND2X1 U1478 ( .A(n1558), .B(n1215), .C(n1214), .D(n1557), .Z(n933) );
  CENXL U1479 ( .A(n1876), .B(n1857), .Z(n1168) );
  CENXL U1480 ( .A(n1857), .B(n1809), .Z(n1163) );
  CENXL U1481 ( .A(n1857), .B(n1810), .Z(n1162) );
  CND2IXL U1482 ( .B(n1876), .A(n1857), .Z(n1169) );
  CIVXL U1483 ( .A(n1834), .Z(n1597) );
  CIVXL U1484 ( .A(n942), .Z(n1598) );
  CIVXL U1485 ( .A(n1598), .Z(n1599) );
  CEN3X2 U1486 ( .A(n1598), .B(n988), .C(n1014), .Z(n670) );
  COND2X1 U1487 ( .A(n1572), .B(n1134), .C(n1133), .D(n1651), .Z(n857) );
  CNIVX4 U1488 ( .A(n1394), .Z(n1818) );
  CNR2X2 U1489 ( .A(n720), .B(n731), .Z(n275) );
  COND2XL U1490 ( .A(n102), .B(n1108), .C(n1107), .D(n100), .Z(n833) );
  CFA1XL U1491 ( .A(n884), .B(n1068), .CI(n960), .CO(n599), .S(n600) );
  CENX2 U1492 ( .A(n1852), .B(a[16]), .Z(n74) );
  CENX1 U1493 ( .A(a[14]), .B(n1855), .Z(n1702) );
  COND2X1 U1494 ( .A(n69), .B(n1184), .C(n1183), .D(n1777), .Z(n904) );
  CND2X2 U1495 ( .A(n1693), .B(n1694), .Z(n888) );
  CND2X2 U1496 ( .A(n1423), .B(n24), .Z(n27) );
  CENXL U1497 ( .A(n1826), .B(n1386), .Z(n1289) );
  CEOX2 U1498 ( .A(n1665), .B(n460), .Z(n450) );
  CENXL U1499 ( .A(n1823), .B(n1390), .Z(n1324) );
  CENXL U1500 ( .A(n1820), .B(b[28]), .Z(n1315) );
  CENXL U1501 ( .A(n1820), .B(b[26]), .Z(n1317) );
  CENXL U1502 ( .A(n1823), .B(b[27]), .Z(n1316) );
  COND2XL U1503 ( .A(n18), .B(n1325), .C(n1324), .D(n1573), .Z(n1039) );
  CIVX2 U1504 ( .A(n1861), .Z(n1857) );
  COND2XL U1505 ( .A(n1653), .B(n1247), .C(n1246), .D(n1576), .Z(n964) );
  COND2XL U1506 ( .A(n1653), .B(n1254), .C(n1253), .D(n1576), .Z(n971) );
  COND2XL U1507 ( .A(n1654), .B(n1236), .C(n1235), .D(n1576), .Z(n953) );
  COND2XL U1508 ( .A(n1654), .B(n1242), .C(n1241), .D(n1576), .Z(n959) );
  COND2XL U1509 ( .A(n1654), .B(n1235), .C(n1234), .D(n1576), .Z(n952) );
  COND2XL U1510 ( .A(n1653), .B(n1234), .C(n1233), .D(n1576), .Z(n951) );
  CENXL U1511 ( .A(n1851), .B(n1813), .Z(n1198) );
  CENXL U1512 ( .A(n1851), .B(n1814), .Z(n1197) );
  CENXL U1513 ( .A(n1851), .B(n1809), .Z(n1203) );
  CENXL U1514 ( .A(n1851), .B(n1815), .Z(n1196) );
  CENXL U1515 ( .A(n1851), .B(n1401), .Z(n1200) );
  CENXL U1516 ( .A(n1851), .B(n1810), .Z(n1202) );
  CENXL U1517 ( .A(n1851), .B(n1805), .Z(n1207) );
  CENXL U1518 ( .A(n1851), .B(n1811), .Z(n1201) );
  CENXL U1519 ( .A(n1851), .B(n1806), .Z(n1206) );
  CENXL U1520 ( .A(n1851), .B(n1807), .Z(n1205) );
  CNIVX4 U1521 ( .A(n1399), .Z(n1813) );
  CENXL U1522 ( .A(n1585), .B(n1817), .Z(n1269) );
  CENXL U1523 ( .A(n1585), .B(n1818), .Z(n1268) );
  CENXL U1524 ( .A(n1585), .B(n1393), .Z(n1267) );
  CENXL U1525 ( .A(n1585), .B(n1816), .Z(n1270) );
  CENXL U1526 ( .A(n1585), .B(n1390), .Z(n1264) );
  CENXL U1527 ( .A(n1836), .B(b[24]), .Z(n1259) );
  CENXL U1528 ( .A(n1833), .B(n1386), .Z(n1260) );
  CENX1 U1529 ( .A(n1780), .B(n1812), .Z(n1159) );
  CIVX3 U1530 ( .A(n1779), .Z(n1780) );
  COND2XL U1531 ( .A(n18), .B(n1315), .C(n1314), .D(n1573), .Z(n1029) );
  COND2XL U1532 ( .A(n18), .B(n1341), .C(n1340), .D(n1573), .Z(n1055) );
  COND2XL U1533 ( .A(n18), .B(n1316), .C(n1315), .D(n1574), .Z(n1030) );
  COND2XL U1534 ( .A(n18), .B(n1336), .C(n1335), .D(n1573), .Z(n1050) );
  COND2XL U1535 ( .A(n18), .B(n1339), .C(n1338), .D(n1574), .Z(n1053) );
  COND2XL U1536 ( .A(n18), .B(n1338), .C(n1337), .D(n1574), .Z(n1052) );
  COND2XL U1537 ( .A(n18), .B(n1326), .C(n1325), .D(n1574), .Z(n1040) );
  COND2XL U1538 ( .A(n18), .B(n1343), .C(n1342), .D(n1573), .Z(n1057) );
  COND2XL U1539 ( .A(n18), .B(n1323), .C(n1322), .D(n1573), .Z(n1037) );
  CIVX2 U1540 ( .A(n1584), .Z(n1833) );
  CIVX2 U1541 ( .A(n1584), .Z(n1836) );
  CEO3XL U1542 ( .A(n699), .B(n701), .C(n703), .Z(n682) );
  CNIVX3 U1543 ( .A(n66), .Z(n1777) );
  CNIVX1 U1544 ( .A(n932), .Z(n1600) );
  COND2XL U1545 ( .A(n61), .B(n1192), .C(n1191), .D(n58), .Z(n911) );
  CENX2 U1546 ( .A(n1835), .B(a[8]), .Z(n42) );
  COND2XL U1547 ( .A(n1559), .B(n1214), .C(n1213), .D(n50), .Z(n932) );
  CENXL U1548 ( .A(n1876), .B(n1828), .Z(n1312) );
  CENXL U1549 ( .A(n1828), .B(n1809), .Z(n1307) );
  CENXL U1550 ( .A(n1828), .B(n1387), .Z(n1290) );
  CENXL U1551 ( .A(n1828), .B(n1806), .Z(n1310) );
  CNIVX4 U1552 ( .A(n1398), .Z(n1814) );
  CENX1 U1553 ( .A(n1843), .B(n1808), .Z(n1252) );
  CNIVX4 U1554 ( .A(n1405), .Z(n1808) );
  CENXL U1555 ( .A(n1857), .B(n1808), .Z(n1164) );
  CENXL U1556 ( .A(n1820), .B(n1808), .Z(n1339) );
  CENXL U1557 ( .A(n1868), .B(n1808), .Z(n1132) );
  CENXL U1558 ( .A(n1831), .B(n1808), .Z(n1308) );
  CENXL U1559 ( .A(n1851), .B(n1808), .Z(n1204) );
  CENXL U1560 ( .A(n1834), .B(n1808), .Z(n1279) );
  CENXL U1561 ( .A(n1862), .B(n1808), .Z(n1147) );
  CNIVX4 U1562 ( .A(n1400), .Z(n1812) );
  COND2X1 U1563 ( .A(n69), .B(n1179), .C(n1178), .D(n1777), .Z(n899) );
  CND2XL U1564 ( .A(n452), .B(n475), .Z(n1635) );
  CEOX1 U1565 ( .A(n452), .B(n475), .Z(n1631) );
  CANR1X1 U1566 ( .A(n301), .B(n1709), .C(n296), .Z(n294) );
  CNIVX2 U1567 ( .A(n900), .Z(n1601) );
  CIVX4 U1568 ( .A(n1846), .Z(n1840) );
  CENXL U1569 ( .A(n1819), .B(n1393), .Z(n1327) );
  CFA1XL U1570 ( .A(n1039), .B(n919), .CI(n961), .CO(n615), .S(n616) );
  CENXL U1571 ( .A(n1828), .B(b[25]), .Z(n1287) );
  CND2X2 U1572 ( .A(n584), .B(n603), .Z(net179871) );
  COR2X1 U1573 ( .A(n583), .B(n562), .Z(net178515) );
  CND2X1 U1574 ( .A(n562), .B(n583), .Z(n212) );
  CND2X1 U1575 ( .A(n604), .B(n623), .Z(n226) );
  CNR2X1 U1576 ( .A(n604), .B(n623), .Z(n225) );
  CFA1X1 U1577 ( .A(net171535), .B(net171537), .CI(net171536), .S(net179596)
         );
  CND2X2 U1578 ( .A(net180046), .B(net180047), .Z(product[27]) );
  CND2X2 U1579 ( .A(net180044), .B(net180045), .Z(net180047) );
  CIVX2 U1580 ( .A(net179917), .Z(net180045) );
  CIVX2 U1581 ( .A(n180), .Z(net180044) );
  CND2X1 U1582 ( .A(n180), .B(net179917), .Z(net180046) );
  CAN2XL U1583 ( .A(n341), .B(n179), .Z(net179917) );
  CIVX2 U1584 ( .A(n176), .Z(n341) );
  CANR1X2 U1585 ( .A(n181), .B(n194), .C(n182), .Z(n180) );
  CIVX2 U1586 ( .A(n195), .Z(n194) );
  CANR1X1 U1587 ( .A(n174), .B(n194), .C(n175), .Z(n173) );
  CENX1 U1588 ( .A(n125), .B(n194), .Z(product[25]) );
  CANR1X1 U1589 ( .A(n196), .B(net179550), .C(n197), .Z(n195) );
  COND1XL U1590 ( .A(n176), .B(n184), .C(n179), .Z(n175) );
  CNR2IXL U1591 ( .B(n181), .A(n176), .Z(n174) );
  CNR2X1 U1592 ( .A(n171), .B(n176), .Z(n169) );
  CND2X1 U1593 ( .A(n169), .B(n181), .Z(n167) );
  CIVX2 U1594 ( .A(n182), .Z(n184) );
  CANR1X1 U1595 ( .A(n196), .B(net179550), .C(n1547), .Z(net181713) );
  CANR1X2 U1596 ( .A(n210), .B(net178516), .C(n201), .Z(n199) );
  CIVX2 U1597 ( .A(n203), .Z(n201) );
  CIVX1 U1598 ( .A(n212), .Z(n210) );
  CIVXL U1599 ( .A(n210), .Z(net179703) );
  CND2X1 U1600 ( .A(net178515), .B(net178516), .Z(n198) );
  CNR2X1 U1601 ( .A(n214), .B(n1578), .Z(n196) );
  CIVXL U1602 ( .A(net179873), .Z(net179908) );
  CIVX2 U1603 ( .A(n222), .Z(n346) );
  CAN2XL U1604 ( .A(n1550), .B(net179908), .Z(net180181) );
  CND2X1 U1605 ( .A(n346), .B(n347), .Z(n214) );
  CIVX2 U1606 ( .A(n226), .Z(n228) );
  CNIVXL U1607 ( .A(n228), .Z(net182652) );
  COR2X1 U1608 ( .A(n540), .B(n561), .Z(net178516) );
  CND2XL U1609 ( .A(net178516), .B(n203), .Z(n126) );
  CND2X1 U1610 ( .A(n561), .B(n540), .Z(n203) );
  CNIVXL U1611 ( .A(net178515), .Z(net180512) );
  CND2XL U1612 ( .A(n226), .B(n347), .Z(n129) );
  CNR2X1 U1613 ( .A(n187), .B(n192), .Z(n181) );
  COND1X2 U1614 ( .A(n193), .B(n187), .C(n188), .Z(n182) );
  COND1XL U1615 ( .A(n233), .B(n245), .C(n234), .Z(net179550) );
  CIVX2 U1616 ( .A(n187), .Z(n342) );
  CIVX2 U1617 ( .A(n192), .Z(n343) );
  COND1X1 U1618 ( .A(n192), .B(net181713), .C(n193), .Z(net178945) );
  CND2XL U1619 ( .A(n343), .B(n193), .Z(n125) );
  CND2XL U1620 ( .A(n342), .B(n188), .Z(n124) );
  CIVXL U1621 ( .A(n214), .Z(n216) );
  CNIVXL U1622 ( .A(n214), .Z(net180533) );
  COAN1X2 U1623 ( .A(n233), .B(n245), .C(n234), .Z(net180264) );
  CIVX2 U1624 ( .A(n245), .Z(n244) );
  COAN1X1 U1625 ( .A(n242), .B(n245), .C(n243), .Z(n239) );
  CNR2X2 U1626 ( .A(n1672), .B(net182652), .Z(n1673) );
  COND2XL U1627 ( .A(n69), .B(n1171), .C(n1170), .D(n1776), .Z(n891) );
  COND2XL U1628 ( .A(n69), .B(n1172), .C(n1171), .D(n1777), .Z(n892) );
  COND2XL U1629 ( .A(n69), .B(n1182), .C(n1181), .D(n1776), .Z(n902) );
  COND2XL U1630 ( .A(n69), .B(n1183), .C(n1182), .D(n1776), .Z(n903) );
  COND2XL U1631 ( .A(n69), .B(n1180), .C(n1179), .D(n1777), .Z(n900) );
  COND2XL U1632 ( .A(n69), .B(n1186), .C(n1185), .D(n1777), .Z(n906) );
  COND2X1 U1633 ( .A(n69), .B(n1187), .C(n1186), .D(n1777), .Z(n907) );
  CENXL U1634 ( .A(n1855), .B(n1818), .Z(n1172) );
  CENXL U1635 ( .A(n1783), .B(n1812), .Z(n1114) );
  CENXL U1636 ( .A(n1841), .B(n1812), .Z(n1247) );
  CENXL U1637 ( .A(n1826), .B(n1812), .Z(n1303) );
  CENXL U1638 ( .A(n1853), .B(n1812), .Z(n1178) );
  CENXL U1639 ( .A(n1864), .B(n1812), .Z(n1142) );
  CENXL U1640 ( .A(n1851), .B(n1812), .Z(n1199) );
  COND1XL U1641 ( .A(n266), .B(n283), .C(n267), .Z(n1602) );
  COND1X1 U1642 ( .A(n266), .B(n283), .C(n267), .Z(n265) );
  COND2X1 U1643 ( .A(n1653), .B(n1250), .C(n1249), .D(n1576), .Z(n967) );
  CNIVX4 U1644 ( .A(n1402), .Z(n1811) );
  CAOR1X1 U1645 ( .A(n1763), .B(n1754), .C(n1757), .Z(n1603) );
  CND2X4 U1646 ( .A(n1417), .B(n74), .Z(n77) );
  CEOX2 U1647 ( .A(n1857), .B(a[16]), .Z(n1417) );
  CND2XL U1648 ( .A(n703), .B(n701), .Z(n1649) );
  CND2X4 U1649 ( .A(n1676), .B(n1677), .Z(product[11]) );
  CEOX2 U1650 ( .A(n538), .B(n559), .Z(n1604) );
  CEOX1 U1651 ( .A(n1604), .B(n557), .Z(n528) );
  CND2XL U1652 ( .A(n557), .B(n559), .Z(n1605) );
  CND2XL U1653 ( .A(n557), .B(n538), .Z(n1606) );
  CND2XL U1654 ( .A(n559), .B(n538), .Z(n1607) );
  CND3X1 U1655 ( .A(n1605), .B(n1606), .C(n1607), .Z(n527) );
  CEO3X2 U1656 ( .A(n868), .B(n1066), .C(n916), .Z(n558) );
  CND2XL U1657 ( .A(n868), .B(n916), .Z(n1608) );
  CND2XL U1658 ( .A(n868), .B(n1066), .Z(n1609) );
  CND2XL U1659 ( .A(n916), .B(n1066), .Z(n1610) );
  CND3X1 U1660 ( .A(n1608), .B(n1609), .C(n1610), .Z(n557) );
  CENXL U1661 ( .A(n1820), .B(n1391), .Z(n1325) );
  CENXL U1662 ( .A(n1822), .B(n1401), .Z(n1335) );
  CENXL U1663 ( .A(n1824), .B(n1812), .Z(n1334) );
  CENXL U1664 ( .A(n1823), .B(n1813), .Z(n1333) );
  COND2X1 U1665 ( .A(n44), .B(n1238), .C(n1237), .D(n1576), .Z(n955) );
  CIVX3 U1666 ( .A(n63), .Z(n1856) );
  CIVX4 U1667 ( .A(n1856), .Z(n1852) );
  COND1X2 U1668 ( .A(n248), .B(n252), .C(n249), .Z(n247) );
  CANR1X4 U1669 ( .A(n1766), .B(n1567), .C(n1753), .Z(n272) );
  CIVX2 U1670 ( .A(n71), .Z(n1861) );
  CEO3X2 U1671 ( .A(n863), .B(n1061), .C(n1617), .Z(n432) );
  CND2XL U1672 ( .A(n863), .B(n1061), .Z(n1611) );
  CND2XL U1673 ( .A(n863), .B(n893), .Z(n1612) );
  CND2XL U1674 ( .A(n1061), .B(n893), .Z(n1613) );
  CND3X1 U1675 ( .A(n1611), .B(n1612), .C(n1613), .Z(n431) );
  CND2X1 U1676 ( .A(n430), .B(n434), .Z(n1614) );
  CND2X1 U1677 ( .A(n430), .B(n432), .Z(n1615) );
  CND2X1 U1678 ( .A(n434), .B(n432), .Z(n1616) );
  CND3X2 U1679 ( .A(n1614), .B(n1615), .C(n1616), .Z(n421) );
  CNIVX1 U1680 ( .A(n893), .Z(n1617) );
  COND2XL U1681 ( .A(n69), .B(n1173), .C(n1172), .D(n1777), .Z(n893) );
  CENX2 U1682 ( .A(n1762), .B(n1618), .Z(product[12]) );
  COND1X1 U1683 ( .A(n1761), .B(n291), .C(n1760), .Z(n1618) );
  CND2X4 U1684 ( .A(n1423), .B(n24), .Z(n1619) );
  CND2X2 U1685 ( .A(n1423), .B(n24), .Z(n1620) );
  CIVX4 U1686 ( .A(n1871), .Z(n1868) );
  CIVXL U1687 ( .A(n864), .Z(n1622) );
  CIVXL U1688 ( .A(n1622), .Z(n1623) );
  CENX2 U1689 ( .A(n257), .B(n133), .Z(product[17]) );
  CFA1X1 U1690 ( .A(n842), .B(n1600), .CI(n852), .CO(n461), .S(n462) );
  CENX1 U1691 ( .A(n1870), .B(n1401), .Z(n1128) );
  CENXL U1692 ( .A(n1583), .B(n1390), .Z(n1189) );
  CENXL U1693 ( .A(n1583), .B(n1391), .Z(n1190) );
  CENXL U1694 ( .A(n1583), .B(n1816), .Z(n1195) );
  CENXL U1695 ( .A(n1583), .B(n1393), .Z(n1192) );
  CENXL U1696 ( .A(n1583), .B(n1817), .Z(n1194) );
  CEOX4 U1697 ( .A(n1756), .B(n1759), .Z(product[10]) );
  CND2X2 U1698 ( .A(n1580), .B(n1675), .Z(n1676) );
  CIVX1 U1699 ( .A(n1768), .Z(n261) );
  CND2X2 U1700 ( .A(n1674), .B(n291), .Z(n1677) );
  CENX1 U1701 ( .A(n127), .B(n213), .Z(product[23]) );
  CFA1X1 U1702 ( .A(n908), .B(n926), .CI(n946), .CO(n729), .S(n730) );
  COND2X1 U1703 ( .A(n97), .B(n1120), .C(n1119), .D(n95), .Z(n844) );
  CNIVX4 U1704 ( .A(n116), .Z(n1875) );
  CND2XL U1705 ( .A(n1599), .B(n1014), .Z(n1626) );
  CND2XL U1706 ( .A(n1599), .B(n988), .Z(n1627) );
  CND2X1 U1707 ( .A(n1014), .B(n988), .Z(n1628) );
  CND3X1 U1708 ( .A(n1626), .B(n1627), .C(n1628), .Z(n669) );
  COND2X1 U1709 ( .A(n61), .B(n1208), .C(n1207), .D(n58), .Z(n927) );
  CENXL U1710 ( .A(n1876), .B(n1583), .Z(n1208) );
  CANR1X2 U1711 ( .A(n1763), .B(n1754), .C(n1757), .Z(n1679) );
  CIVXL U1712 ( .A(n104), .Z(n1437) );
  CENXL U1713 ( .A(n1808), .B(n104), .Z(n1099) );
  CENXL U1714 ( .A(n1806), .B(n104), .Z(n1101) );
  CENXL U1715 ( .A(n1807), .B(n104), .Z(n1100) );
  CENXL U1716 ( .A(n1809), .B(n1593), .Z(n1098) );
  COND2X1 U1717 ( .A(n36), .B(n1273), .C(n1272), .D(n1796), .Z(n989) );
  CENXL U1718 ( .A(n1820), .B(n1387), .Z(n1321) );
  CENXL U1719 ( .A(n1839), .B(n1387), .Z(n1234) );
  CENXL U1720 ( .A(n1836), .B(n1387), .Z(n1261) );
  CNIVX4 U1721 ( .A(n66), .Z(n1775) );
  CENX2 U1722 ( .A(n1851), .B(a[14]), .Z(n66) );
  CND2X2 U1723 ( .A(n1412), .B(n105), .Z(n107) );
  CIVX1 U1724 ( .A(n1018), .Z(n1629) );
  CIVX2 U1725 ( .A(n1629), .Z(n1630) );
  CEO3X2 U1726 ( .A(n489), .B(n485), .C(n487), .Z(n454) );
  CND2X1 U1727 ( .A(n489), .B(n487), .Z(n1633) );
  CND3X2 U1728 ( .A(n1632), .B(n1633), .C(n1634), .Z(n453) );
  CND2X1 U1729 ( .A(n475), .B(n454), .Z(n1637) );
  CND3X1 U1730 ( .A(n1635), .B(n1636), .C(n1637), .Z(n445) );
  CIVX2 U1731 ( .A(n165), .Z(n163) );
  CANR1XL U1732 ( .A(n163), .B(net178510), .C(n158), .Z(n156) );
  COR2X1 U1733 ( .A(n412), .B(n439), .Z(net178506) );
  CND2XL U1734 ( .A(net178506), .B(n165), .Z(net178944) );
  CND2X1 U1735 ( .A(n412), .B(n439), .Z(n165) );
  COND1X1 U1736 ( .A(n167), .B(net181713), .C(n168), .Z(net182753) );
  CIVXL U1737 ( .A(n171), .Z(n340) );
  CND2XL U1738 ( .A(n340), .B(n172), .Z(n122) );
  COR2X1 U1739 ( .A(n384), .B(n411), .Z(net178510) );
  CND2X1 U1740 ( .A(n384), .B(n411), .Z(n160) );
  CIVXL U1741 ( .A(n160), .Z(n158) );
  CHA1X1 U1742 ( .A(n811), .B(n1045), .CO(n717), .S(n718) );
  COND2X1 U1743 ( .A(n69), .B(n1856), .C(n1188), .D(n1777), .Z(n811) );
  CEOX2 U1744 ( .A(a[2]), .B(n1821), .Z(n1424) );
  CENX2 U1745 ( .A(n1852), .B(a[16]), .Z(n1638) );
  CENX2 U1746 ( .A(n1852), .B(a[16]), .Z(n1639) );
  COND2X1 U1747 ( .A(n1570), .B(n1277), .C(n1276), .D(n1796), .Z(n993) );
  CENXL U1748 ( .A(n1861), .B(a[18]), .Z(n1704) );
  CIVX1 U1749 ( .A(n291), .Z(n1675) );
  CENXL U1750 ( .A(n1807), .B(n109), .Z(n1093) );
  CND2IXL U1751 ( .B(n1876), .A(n109), .Z(n1097) );
  CENXL U1752 ( .A(n109), .B(a[30]), .Z(n114) );
  CENXL U1753 ( .A(n1805), .B(n109), .Z(n1095) );
  CENXL U1754 ( .A(n1806), .B(n109), .Z(n1094) );
  CEOX2 U1755 ( .A(a[28]), .B(n109), .Z(n1411) );
  COND2XL U1756 ( .A(n61), .B(n1201), .C(n1200), .D(n58), .Z(n920) );
  COND2XL U1757 ( .A(n61), .B(n1200), .C(n1199), .D(n58), .Z(n919) );
  COND2XL U1758 ( .A(n61), .B(n1197), .C(n1196), .D(n58), .Z(n916) );
  CENXL U1759 ( .A(n1849), .B(n1808), .Z(n1227) );
  CENXL U1760 ( .A(n1864), .B(n1813), .Z(n1141) );
  CENXL U1761 ( .A(n1864), .B(n1814), .Z(n1140) );
  CENXL U1762 ( .A(n1864), .B(n1401), .Z(n1143) );
  CIVX2 U1763 ( .A(n79), .Z(n1867) );
  CIVX1 U1764 ( .A(n1847), .Z(n1842) );
  CEO3X2 U1765 ( .A(n684), .B(n695), .C(n682), .Z(n678) );
  CEOX2 U1766 ( .A(n680), .B(n693), .Z(n1640) );
  CEOX2 U1767 ( .A(n1640), .B(n678), .Z(n676) );
  CND2XL U1768 ( .A(n684), .B(n695), .Z(n1641) );
  CND2XL U1769 ( .A(n684), .B(n682), .Z(n1642) );
  CND2XL U1770 ( .A(n695), .B(n682), .Z(n1643) );
  CND3X1 U1771 ( .A(n1641), .B(n1642), .C(n1643), .Z(n677) );
  CND2XL U1772 ( .A(n680), .B(n693), .Z(n1644) );
  CND2XL U1773 ( .A(n680), .B(n678), .Z(n1645) );
  CND2XL U1774 ( .A(n693), .B(n678), .Z(n1646) );
  CND3XL U1775 ( .A(n1644), .B(n1645), .C(n1646), .Z(n675) );
  CND2XL U1776 ( .A(n699), .B(n703), .Z(n1647) );
  CND2XL U1777 ( .A(n699), .B(n701), .Z(n1648) );
  CND3X1 U1778 ( .A(n1647), .B(n1648), .C(n1649), .Z(n681) );
  CAN2X2 U1779 ( .A(n1772), .B(n1767), .Z(n1700) );
  CENXL U1780 ( .A(n1805), .B(n104), .Z(n1102) );
  CENX1 U1781 ( .A(n1805), .B(n1873), .Z(n1111) );
  CENX1 U1782 ( .A(n1862), .B(a[20]), .Z(n1650) );
  CENX1 U1783 ( .A(n1862), .B(a[20]), .Z(n1651) );
  COND2X1 U1784 ( .A(n1571), .B(n1276), .C(n1275), .D(n1796), .Z(n992) );
  CENX1 U1785 ( .A(n1588), .B(n1814), .Z(n1301) );
  CNIVX2 U1786 ( .A(n1696), .Z(n1652) );
  CENXL U1787 ( .A(n1853), .B(n1401), .Z(n1179) );
  CENXL U1788 ( .A(n1854), .B(n1807), .Z(n1184) );
  CENXL U1789 ( .A(n1854), .B(n1806), .Z(n1185) );
  CENXL U1790 ( .A(n1854), .B(n1805), .Z(n1186) );
  CND2X4 U1791 ( .A(n1421), .B(n1576), .Z(n1654) );
  CND2X1 U1792 ( .A(n1421), .B(n1575), .Z(n44) );
  CEOX2 U1793 ( .A(a[8]), .B(n1844), .Z(n1421) );
  CND2X2 U1794 ( .A(n129), .B(net180393), .Z(n1655) );
  CND2X2 U1795 ( .A(n1655), .B(n1656), .Z(product[21]) );
  CIVX2 U1796 ( .A(n86), .Z(n1871) );
  COND2XL U1797 ( .A(n18), .B(n1329), .C(n1328), .D(n1573), .Z(n1043) );
  CIVX2 U1798 ( .A(n99), .Z(n1874) );
  CND2XL U1799 ( .A(n1873), .B(n1809), .Z(n1659) );
  CND2X2 U1800 ( .A(n1657), .B(n1658), .Z(n1660) );
  CND2X2 U1801 ( .A(n1659), .B(n1660), .Z(n1107) );
  CIVXL U1802 ( .A(n1873), .Z(n1657) );
  CIVX1 U1803 ( .A(n1809), .Z(n1658) );
  CNIVX4 U1804 ( .A(n1404), .Z(n1809) );
  CND2IXL U1805 ( .B(n1876), .A(n113), .Z(n1092) );
  CENXL U1806 ( .A(n1805), .B(n113), .Z(n1090) );
  CENXL U1807 ( .A(n1841), .B(n1401), .Z(n1248) );
  CENXL U1808 ( .A(n1841), .B(n1815), .Z(n1244) );
  CNR2XL U1809 ( .A(n1248), .B(n1575), .Z(n1717) );
  CENXL U1810 ( .A(n1841), .B(n1386), .Z(n1233) );
  COND2X1 U1811 ( .A(n1572), .B(n1129), .C(n1128), .D(n1650), .Z(n852) );
  CIVXL U1812 ( .A(n86), .Z(n1872) );
  CENX2 U1813 ( .A(n272), .B(n1700), .Z(product[15]) );
  CIVX2 U1814 ( .A(n1754), .Z(n291) );
  CND2X1 U1815 ( .A(n1591), .B(net180393), .Z(n1661) );
  CND2X1 U1816 ( .A(n1661), .B(n206), .Z(n204) );
  CENXL U1817 ( .A(n1849), .B(n1813), .Z(n1221) );
  CENXL U1818 ( .A(n1849), .B(n1814), .Z(n1220) );
  CENXL U1819 ( .A(n1849), .B(n1812), .Z(n1222) );
  CENXL U1820 ( .A(n1849), .B(n1815), .Z(n1219) );
  CENXL U1821 ( .A(n1849), .B(n1817), .Z(n1217) );
  CENXL U1822 ( .A(n1849), .B(n1393), .Z(n1215) );
  CENXL U1823 ( .A(n1849), .B(n1818), .Z(n1216) );
  CENXL U1824 ( .A(n1849), .B(n1391), .Z(n1213) );
  CENXL U1825 ( .A(n1826), .B(n1815), .Z(n1300) );
  CENXL U1826 ( .A(n1588), .B(n1816), .Z(n1299) );
  CENXL U1827 ( .A(n1827), .B(n1817), .Z(n1298) );
  CEOX2 U1828 ( .A(a[6]), .B(n1837), .Z(n1422) );
  COND2XL U1829 ( .A(n107), .B(n1099), .C(n1098), .D(n105), .Z(n825) );
  COND2XL U1830 ( .A(n107), .B(n1101), .C(n1100), .D(n105), .Z(n827) );
  CENXL U1831 ( .A(n1873), .B(n1811), .Z(n1105) );
  CND2IXL U1832 ( .B(n1876), .A(n1873), .Z(n1113) );
  CENXL U1833 ( .A(n1873), .B(n1810), .Z(n1106) );
  CENXL U1834 ( .A(n1873), .B(n1806), .Z(n1110) );
  CEO3X1 U1835 ( .A(n486), .B(n488), .C(n505), .Z(n476) );
  CND2XL U1836 ( .A(n486), .B(n505), .Z(n1662) );
  CND2XL U1837 ( .A(n486), .B(n488), .Z(n1663) );
  CND2X1 U1838 ( .A(n505), .B(n488), .Z(n1664) );
  CND3X1 U1839 ( .A(n1662), .B(n1663), .C(n1664), .Z(n475) );
  CFA1X1 U1840 ( .A(n994), .B(n1078), .CI(n1048), .CO(n749), .S(n750) );
  COND2X1 U1841 ( .A(n1571), .B(n1278), .C(n1277), .D(n1796), .Z(n994) );
  CND2X2 U1842 ( .A(n110), .B(n1411), .Z(n112) );
  COND1X1 U1843 ( .A(n251), .B(n264), .C(n252), .Z(n250) );
  CENX2 U1844 ( .A(n250), .B(n132), .Z(product[18]) );
  CENXL U1845 ( .A(n1875), .B(n113), .Z(n1091) );
  CENXL U1846 ( .A(n1875), .B(n1824), .Z(n1343) );
  CENXL U1847 ( .A(n1875), .B(n1783), .Z(n1123) );
  CENXL U1848 ( .A(n1875), .B(n1837), .Z(n1283) );
  CENXL U1849 ( .A(n1875), .B(n1870), .Z(n1136) );
  CENXL U1850 ( .A(n1875), .B(n1844), .Z(n1256) );
  CENXL U1851 ( .A(n1875), .B(n109), .Z(n1096) );
  CENXL U1852 ( .A(n1875), .B(n1855), .Z(n1187) );
  CENXL U1853 ( .A(n1875), .B(n1865), .Z(n1151) );
  CENXL U1854 ( .A(n1875), .B(n1593), .Z(n1103) );
  CNIVX4 U1855 ( .A(n1406), .Z(n1807) );
  CIVX2 U1856 ( .A(n1683), .Z(n348) );
  CNR2X1 U1857 ( .A(n1549), .B(net180090), .Z(n1672) );
  COND2X1 U1858 ( .A(n1570), .B(n1272), .C(n1271), .D(n1796), .Z(n988) );
  CND2IXL U1859 ( .B(n275), .A(n276), .Z(n136) );
  COND2X1 U1860 ( .A(n1558), .B(n1230), .C(n1229), .D(n50), .Z(n948) );
  COND2X1 U1861 ( .A(n53), .B(n1228), .C(n1227), .D(n50), .Z(n946) );
  CIVX8 U1862 ( .A(n1798), .Z(n24) );
  CND2X4 U1863 ( .A(n1794), .B(n1795), .Z(n1798) );
  CIVX2 U1864 ( .A(n1825), .Z(n1821) );
  CND2IX4 U1865 ( .B(n1702), .A(n1775), .Z(n69) );
  CEO3X2 U1866 ( .A(n864), .B(n1062), .C(n912), .Z(n460) );
  CEOX2 U1867 ( .A(n462), .B(n456), .Z(n1665) );
  CND2XL U1868 ( .A(n1623), .B(n1062), .Z(n1666) );
  CND2XL U1869 ( .A(n1623), .B(n912), .Z(n1667) );
  CND2XL U1870 ( .A(n1062), .B(n912), .Z(n1668) );
  CND2XL U1871 ( .A(n462), .B(n456), .Z(n1669) );
  CND2XL U1872 ( .A(n462), .B(n460), .Z(n1670) );
  CND2XL U1873 ( .A(n456), .B(n460), .Z(n1671) );
  CND3X1 U1874 ( .A(n1669), .B(n1670), .C(n1671), .Z(n449) );
  CIVX2 U1875 ( .A(n139), .Z(n1674) );
  CEOX2 U1876 ( .A(a[24]), .B(n1873), .Z(n1413) );
  CENXL U1877 ( .A(n1849), .B(n1388), .Z(n1210) );
  CENXL U1878 ( .A(n1849), .B(n1389), .Z(n1211) );
  CENXL U1879 ( .A(n1849), .B(n1816), .Z(n1218) );
  CENXL U1880 ( .A(n1849), .B(n1811), .Z(n1224) );
  CENXL U1881 ( .A(n1849), .B(n1809), .Z(n1226) );
  CENXL U1882 ( .A(n1849), .B(n1401), .Z(n1223) );
  CENXL U1883 ( .A(n1849), .B(n1810), .Z(n1225) );
  CENXL U1884 ( .A(n1849), .B(n1807), .Z(n1228) );
  CENXL U1885 ( .A(n1849), .B(n1805), .Z(n1230) );
  CENXL U1886 ( .A(n1849), .B(n1806), .Z(n1229) );
  CENXL U1887 ( .A(n1875), .B(n1873), .Z(n1112) );
  CNR2X2 U1888 ( .A(n732), .B(n743), .Z(n280) );
  CENXL U1889 ( .A(n1875), .B(n1849), .Z(n1231) );
  CIVXL U1890 ( .A(n347), .Z(net180090) );
  CIVX2 U1891 ( .A(n225), .Z(n347) );
  CANR1X1 U1892 ( .A(n1763), .B(n1754), .C(n1757), .Z(n283) );
  CEOX1 U1893 ( .A(n1758), .B(n1732), .Z(n540) );
  CENX1 U1894 ( .A(net178944), .B(net182753), .Z(product[29]) );
  CENX2 U1895 ( .A(n126), .B(n204), .Z(product[24]) );
  CANR1X2 U1896 ( .A(n1771), .B(n1678), .C(n279), .Z(n1701) );
  COND1X1 U1897 ( .A(n1549), .B(net180533), .C(net179577), .Z(n213) );
  COND2X1 U1898 ( .A(n1620), .B(n1293), .C(n1292), .D(n24), .Z(n1008) );
  CENXL U1899 ( .A(n1826), .B(n1389), .Z(n1292) );
  CENXL U1900 ( .A(n1830), .B(n1390), .Z(n1293) );
  CIVX1 U1901 ( .A(n1867), .Z(n1863) );
  CIVXL U1902 ( .A(n1867), .Z(n1864) );
  CENX4 U1903 ( .A(a[10]), .B(n1840), .Z(n50) );
  CNR2IX1 U1904 ( .B(n1876), .A(n50), .Z(n950) );
  CENX4 U1905 ( .A(n1868), .B(a[22]), .Z(n95) );
  CENXL U1906 ( .A(n93), .B(n1807), .Z(n1120) );
  COND2XL U1907 ( .A(n107), .B(n1437), .C(n105), .D(n1104), .Z(n805) );
  CFA1X1 U1908 ( .A(n894), .B(n1004), .CI(n978), .CO(n455), .S(n456) );
  COND2X1 U1909 ( .A(n1570), .B(n1262), .C(n1261), .D(n1796), .Z(n978) );
  CENXL U1910 ( .A(n144), .B(n318), .Z(product[6]) );
  COND1X1 U1911 ( .A(n321), .B(n319), .C(n320), .Z(n318) );
  CANR1X1 U1912 ( .A(n1708), .B(n310), .C(n307), .Z(n305) );
  CEOX1 U1913 ( .A(a[26]), .B(n104), .Z(n1412) );
  CENXL U1914 ( .A(n1824), .B(n1818), .Z(n1328) );
  CENXL U1915 ( .A(n1820), .B(n1815), .Z(n1331) );
  CENXL U1916 ( .A(n1819), .B(n1816), .Z(n1330) );
  CFA1X1 U1917 ( .A(n1072), .B(n922), .CI(n1042), .CO(n671), .S(n672) );
  CIVXL U1918 ( .A(net179703), .Z(net179704) );
  CENXL U1919 ( .A(n1873), .B(n1807), .Z(n1109) );
  CENX2 U1920 ( .A(n1873), .B(a[26]), .Z(n105) );
  CENX4 U1921 ( .A(n1848), .B(a[12]), .Z(n58) );
  CENXL U1922 ( .A(n1583), .B(n1818), .Z(n1193) );
  CND2XL U1923 ( .A(n173), .B(net179450), .Z(n1682) );
  CENX2 U1924 ( .A(n1728), .B(n1680), .Z(n624) );
  CENX2 U1925 ( .A(n1729), .B(n1725), .Z(n1680) );
  CNR2X2 U1926 ( .A(n624), .B(n1727), .Z(n1683) );
  CEOX1 U1927 ( .A(a[22]), .B(n93), .Z(n1414) );
  CND2X4 U1928 ( .A(n1419), .B(n58), .Z(n61) );
  COND2X1 U1929 ( .A(n1558), .B(n1213), .C(n1212), .D(n50), .Z(n931) );
  CENXL U1930 ( .A(n1849), .B(n1390), .Z(n1212) );
  CENXL U1931 ( .A(n1843), .B(n1392), .Z(n1239) );
  CENXL U1932 ( .A(n1819), .B(n1392), .Z(n1326) );
  CENXL U1933 ( .A(n1849), .B(n1392), .Z(n1214) );
  CENXL U1934 ( .A(n1837), .B(n1392), .Z(n1266) );
  CENXL U1935 ( .A(n1855), .B(n1392), .Z(n1170) );
  CENXL U1936 ( .A(n1828), .B(n1392), .Z(n1295) );
  CENXL U1937 ( .A(n1583), .B(n1392), .Z(n1191) );
  CEOX2 U1938 ( .A(n1652), .B(n239), .Z(product[20]) );
  CIVX4 U1939 ( .A(n1874), .Z(n1873) );
  CENX2 U1940 ( .A(n124), .B(net178945), .Z(product[26]) );
  CENX2 U1941 ( .A(n93), .B(a[24]), .Z(n100) );
  COND2X1 U1942 ( .A(n102), .B(n1109), .C(n1108), .D(n100), .Z(n834) );
  CND2X1 U1943 ( .A(n624), .B(n1727), .Z(n238) );
  CND2X2 U1944 ( .A(n1413), .B(n100), .Z(n102) );
  COND2XL U1945 ( .A(n102), .B(n1874), .C(n100), .D(n1113), .Z(n806) );
  COND2XL U1946 ( .A(n102), .B(n1106), .C(n1105), .D(n100), .Z(n831) );
  COND1X2 U1947 ( .A(n1769), .B(n264), .C(n1768), .Z(n257) );
  CND2X1 U1948 ( .A(net179451), .B(n122), .Z(n1681) );
  CND2X2 U1949 ( .A(n1681), .B(n1682), .Z(product[28]) );
  CIVX2 U1950 ( .A(n122), .Z(net179450) );
  CIVXL U1951 ( .A(n173), .Z(net179451) );
  CND2XL U1952 ( .A(n1728), .B(n1725), .Z(n1684) );
  CND2XL U1953 ( .A(n1728), .B(n1729), .Z(n1685) );
  CND2XL U1954 ( .A(n1725), .B(n1729), .Z(n1686) );
  CND3XL U1955 ( .A(n1684), .B(n1685), .C(n1686), .Z(n623) );
  CND2X1 U1956 ( .A(n674), .B(n672), .Z(n1687) );
  CND2X1 U1957 ( .A(n674), .B(n685), .Z(n1688) );
  CND2X1 U1958 ( .A(n672), .B(n685), .Z(n1689) );
  CND3X2 U1959 ( .A(n1687), .B(n1688), .C(n1689), .Z(n665) );
  CENXL U1960 ( .A(n1852), .B(n1810), .Z(n1181) );
  CENXL U1961 ( .A(n1852), .B(n1808), .Z(n1183) );
  CENXL U1962 ( .A(n1852), .B(n1809), .Z(n1182) );
  CIVX1 U1963 ( .A(n1825), .Z(n1824) );
  COR2X1 U1964 ( .A(n329), .B(n327), .Z(n1690) );
  CND2X2 U1965 ( .A(n1690), .B(n328), .Z(n326) );
  CNR2X1 U1966 ( .A(n802), .B(n1087), .Z(n327) );
  CANR1X2 U1967 ( .A(n326), .B(n1710), .C(n323), .Z(n321) );
  CENXL U1968 ( .A(n146), .B(n326), .Z(product[4]) );
  CNR2XL U1969 ( .A(n18), .B(n1342), .Z(n1691) );
  CNR2XL U1970 ( .A(n1341), .B(n1574), .Z(n1692) );
  COR2X1 U1971 ( .A(n1691), .B(n1692), .Z(n1056) );
  CENXL U1972 ( .A(n1822), .B(n1805), .Z(n1342) );
  CENXL U1973 ( .A(n1819), .B(n1806), .Z(n1341) );
  CIVX4 U1974 ( .A(n1582), .Z(n1851) );
  CENX1 U1975 ( .A(n1858), .B(n1806), .Z(n1166) );
  CENX1 U1976 ( .A(n1858), .B(n1805), .Z(n1167) );
  COR2XL U1977 ( .A(n77), .B(n1167), .Z(n1693) );
  COR2XL U1978 ( .A(n1166), .B(n1639), .Z(n1694) );
  CNR2X1 U1979 ( .A(n692), .B(n705), .Z(n258) );
  CND2X1 U1980 ( .A(n754), .B(n763), .Z(n290) );
  COR2X1 U1981 ( .A(n800), .B(n801), .Z(n1710) );
  CNR2IX1 U1982 ( .B(n1876), .A(n1776), .Z(n908) );
  CNR2IX1 U1983 ( .B(n1876), .A(n114), .Z(n820) );
  CNR2IX1 U1984 ( .B(n1876), .A(n1638), .Z(n890) );
  CNR2IX1 U1985 ( .B(n1876), .A(n1781), .Z(n874) );
  CIVX2 U1986 ( .A(n1767), .Z(n269) );
  CENX1 U1987 ( .A(a[18]), .B(n1865), .Z(n1719) );
  CENX1 U1988 ( .A(n1603), .B(n1703), .Z(product[13]) );
  CND2XL U1989 ( .A(n1773), .B(n352), .Z(n251) );
  CND2XL U1990 ( .A(n1709), .B(n1594), .Z(n293) );
  CNR2XL U1991 ( .A(n286), .B(n289), .Z(n284) );
  CND2XL U1992 ( .A(n706), .B(n719), .Z(n271) );
  CND2XL U1993 ( .A(n676), .B(n691), .Z(n256) );
  CND2XL U1994 ( .A(n1709), .B(n298), .Z(n140) );
  CND2IXL U1995 ( .B(n286), .A(n287), .Z(n138) );
  COND1X1 U1996 ( .A(n311), .B(n313), .C(n312), .Z(n310) );
  CND2IXL U1997 ( .B(n311), .A(n312), .Z(n143) );
  CND2XL U1998 ( .A(n363), .B(n320), .Z(n145) );
  CEOXL U1999 ( .A(n321), .B(n145), .Z(product[5]) );
  CND2XL U2000 ( .A(n1712), .B(n317), .Z(n144) );
  CND2XL U2001 ( .A(n744), .B(n753), .Z(n287) );
  CND2XL U2002 ( .A(n1710), .B(n325), .Z(n146) );
  CND3X1 U2003 ( .A(n1789), .B(n1790), .C(n1791), .Z(n699) );
  CEOX1 U2004 ( .A(n1695), .B(n966), .Z(n700) );
  CEOX1 U2005 ( .A(n990), .B(n1016), .Z(n1695) );
  COR2XL U2006 ( .A(n1088), .B(n1058), .Z(n1713) );
  CNIVX4 U2007 ( .A(n33), .Z(n1796) );
  CND2XL U2008 ( .A(n238), .B(n348), .Z(n1696) );
  CIVXL U2009 ( .A(n1846), .Z(n1841) );
  CNR2IXL U2010 ( .B(n1876), .A(n1576), .Z(n974) );
  CNR2IXL U2011 ( .B(n1876), .A(n95), .Z(n848) );
  COND2XL U2012 ( .A(n84), .B(n1148), .C(n1147), .D(n1781), .Z(n870) );
  CNR2IXL U2013 ( .B(n1876), .A(n100), .Z(n838) );
  CNR2X1 U2014 ( .A(n44), .B(n1249), .Z(n1716) );
  CEO3X1 U2015 ( .A(n1697), .B(n1698), .C(n399), .Z(n373) );
  CEO3XL U2016 ( .A(n875), .B(n951), .C(n1029), .Z(n1697) );
  CEO3X1 U2017 ( .A(n929), .B(n975), .C(n1001), .Z(n1698) );
  CNR2IXL U2018 ( .B(n1876), .A(n6), .Z(product[0]) );
  CENX2 U2019 ( .A(n1862), .B(a[20]), .Z(n89) );
  CNIVX2 U2020 ( .A(n1395), .Z(n1817) );
  CNIVX4 U2021 ( .A(n1407), .Z(n1806) );
  COR2X2 U2022 ( .A(n1719), .B(n1704), .Z(n84) );
  CNIVX3 U2023 ( .A(n1403), .Z(n1810) );
  CNIVX4 U2024 ( .A(n1408), .Z(n1805) );
  CND2X1 U2025 ( .A(n1766), .B(n1772), .Z(n266) );
  CND2X2 U2026 ( .A(n1792), .B(a[4]), .Z(n1795) );
  CND2XL U2027 ( .A(n114), .B(n1410), .Z(n115) );
  CND2X1 U2028 ( .A(n1771), .B(n1764), .Z(n1703) );
  CENX1 U2029 ( .A(n1586), .B(n152), .Z(product[31]) );
  CENX1 U2030 ( .A(n141), .B(n304), .Z(product[9]) );
  CND2X1 U2031 ( .A(n1708), .B(n309), .Z(n142) );
  CANR1XL U2032 ( .A(n1594), .B(n304), .C(n301), .Z(n299) );
  COND1XL U2033 ( .A(n281), .B(n275), .C(n276), .Z(n274) );
  COND1XL U2034 ( .A(n290), .B(n286), .C(n287), .Z(n285) );
  CEOX1 U2035 ( .A(n563), .B(n544), .Z(n1799) );
  COND1XL U2036 ( .A(n305), .B(n293), .C(n294), .Z(n292) );
  CNR2XL U2037 ( .A(n275), .B(n280), .Z(n273) );
  CND2X1 U2038 ( .A(n692), .B(n705), .Z(n259) );
  COR2X1 U2039 ( .A(n676), .B(n691), .Z(n1705) );
  COR2X1 U2040 ( .A(n719), .B(n706), .Z(n1706) );
  CNR2X1 U2041 ( .A(n744), .B(n753), .Z(n286) );
  CNR2X1 U2042 ( .A(n754), .B(n763), .Z(n289) );
  COR2X1 U2043 ( .A(n772), .B(n779), .Z(n1707) );
  COR2X1 U2044 ( .A(n780), .B(n785), .Z(n1708) );
  COR2X1 U2045 ( .A(n771), .B(n764), .Z(n1709) );
  CND2X1 U2046 ( .A(n772), .B(n779), .Z(n303) );
  CND2X1 U2047 ( .A(n764), .B(n771), .Z(n298) );
  CND2X1 U2048 ( .A(n780), .B(n785), .Z(n309) );
  CND2X1 U2049 ( .A(n732), .B(n743), .Z(n281) );
  CANR1XL U2050 ( .A(n1592), .B(net182753), .C(n154), .Z(n152) );
  CANR1XL U2051 ( .A(net180512), .B(n1551), .C(net179704), .Z(n206) );
  CNR2X1 U2052 ( .A(n786), .B(n791), .Z(n311) );
  CNR2X1 U2053 ( .A(n796), .B(n799), .Z(n319) );
  CENX1 U2054 ( .A(n902), .B(n1711), .Z(n638) );
  CENX1 U2055 ( .A(n1070), .B(n1012), .Z(n1711) );
  CND2X1 U2056 ( .A(n786), .B(n791), .Z(n312) );
  CND2X1 U2057 ( .A(n796), .B(n799), .Z(n320) );
  CND2XL U2058 ( .A(n802), .B(n1087), .Z(n328) );
  CND2X1 U2059 ( .A(n800), .B(n801), .Z(n325) );
  CND2X1 U2060 ( .A(n792), .B(n795), .Z(n317) );
  CND2X1 U2061 ( .A(n1088), .B(n1058), .Z(n333) );
  COR2X1 U2062 ( .A(n792), .B(n795), .Z(n1712) );
  CIVX2 U2063 ( .A(n1797), .Z(n1834) );
  CIVX2 U2064 ( .A(n1821), .Z(n1792) );
  CNR2X2 U2065 ( .A(n492), .B(n515), .Z(n187) );
  CENX1 U2066 ( .A(n244), .B(n131), .Z(product[19]) );
  CND2XL U2067 ( .A(n349), .B(n243), .Z(n131) );
  CENX1 U2068 ( .A(n1869), .B(n1814), .Z(n1125) );
  CND2XL U2069 ( .A(n350), .B(n249), .Z(n132) );
  CENX1 U2070 ( .A(n1836), .B(n1812), .Z(n1274) );
  CENX1 U2071 ( .A(n1870), .B(n1812), .Z(n1127) );
  CENX1 U2072 ( .A(n1842), .B(n1813), .Z(n1246) );
  CENX1 U2073 ( .A(n1840), .B(n1806), .Z(n1254) );
  CENX1 U2074 ( .A(n1819), .B(n1807), .Z(n1340) );
  CENX1 U2075 ( .A(n1840), .B(n1805), .Z(n1255) );
  CENX1 U2076 ( .A(n1854), .B(n1817), .Z(n1173) );
  CENX1 U2077 ( .A(n1840), .B(n1807), .Z(n1253) );
  CENX1 U2078 ( .A(n1862), .B(n1810), .Z(n1145) );
  CENX1 U2079 ( .A(n1854), .B(n1815), .Z(n1175) );
  CENX1 U2080 ( .A(n1853), .B(n1813), .Z(n1177) );
  CENX1 U2081 ( .A(n1853), .B(n1814), .Z(n1176) );
  CENX1 U2082 ( .A(n1853), .B(n1811), .Z(n1180) );
  CENX1 U2083 ( .A(n1862), .B(n1809), .Z(n1146) );
  CENX1 U2084 ( .A(n1843), .B(n1817), .Z(n1242) );
  CENX1 U2085 ( .A(n1824), .B(n1809), .Z(n1338) );
  CENX1 U2086 ( .A(n1839), .B(n1811), .Z(n1249) );
  CENX1 U2087 ( .A(n1869), .B(n1811), .Z(n1129) );
  CENX1 U2088 ( .A(n1836), .B(n1813), .Z(n1273) );
  CENX1 U2089 ( .A(n1870), .B(n1813), .Z(n1126) );
  CENX1 U2090 ( .A(n1826), .B(n1818), .Z(n1297) );
  CENX1 U2091 ( .A(n1833), .B(n1401), .Z(n1275) );
  CENX1 U2092 ( .A(n1588), .B(n1813), .Z(n1302) );
  CENX1 U2093 ( .A(n1830), .B(n1401), .Z(n1304) );
  CENX1 U2094 ( .A(n1834), .B(n1806), .Z(n1281) );
  CENX1 U2095 ( .A(n1836), .B(n1805), .Z(n1282) );
  CENX1 U2096 ( .A(n1836), .B(n1815), .Z(n1271) );
  CENX1 U2097 ( .A(n1833), .B(n1810), .Z(n1277) );
  CENX1 U2098 ( .A(n1833), .B(n1811), .Z(n1276) );
  CENX1 U2099 ( .A(n1860), .B(n1818), .Z(n1153) );
  CNR2IXL U2100 ( .B(n1876), .A(n1573), .Z(n1058) );
  CENX1 U2101 ( .A(n1869), .B(n1805), .Z(n1135) );
  CENX1 U2102 ( .A(n1863), .B(n1807), .Z(n1148) );
  CENX1 U2103 ( .A(n1783), .B(n1808), .Z(n1119) );
  CENX1 U2104 ( .A(n1780), .B(n1813), .Z(n1158) );
  CENX1 U2105 ( .A(n1783), .B(n1401), .Z(n1115) );
  CENX1 U2106 ( .A(n1858), .B(n1807), .Z(n1165) );
  CENX1 U2107 ( .A(n1858), .B(n1401), .Z(n1160) );
  CENX1 U2108 ( .A(n1783), .B(n1811), .Z(n1116) );
  CENX1 U2109 ( .A(n1842), .B(n1810), .Z(n1250) );
  CENX1 U2110 ( .A(n1783), .B(n1809), .Z(n1118) );
  CENX1 U2111 ( .A(n1783), .B(n1810), .Z(n1117) );
  CENX1 U2112 ( .A(n1860), .B(n1817), .Z(n1154) );
  CENX1 U2113 ( .A(n1783), .B(n1805), .Z(n1122) );
  CENX1 U2114 ( .A(n1827), .B(n1810), .Z(n1306) );
  CENX1 U2115 ( .A(n1844), .B(n1809), .Z(n1251) );
  CENX1 U2116 ( .A(n1863), .B(n1805), .Z(n1150) );
  CENX1 U2117 ( .A(n1865), .B(n1815), .Z(n1139) );
  CENX1 U2118 ( .A(n1780), .B(n1815), .Z(n1156) );
  CENX1 U2119 ( .A(n1843), .B(n1818), .Z(n1241) );
  CENX1 U2120 ( .A(n1820), .B(n1811), .Z(n1336) );
  CENX1 U2121 ( .A(n1863), .B(n1811), .Z(n1144) );
  CENX1 U2122 ( .A(n1824), .B(n1810), .Z(n1337) );
  CENX1 U2123 ( .A(n1826), .B(n1811), .Z(n1305) );
  CENX1 U2124 ( .A(n1869), .B(n1806), .Z(n1134) );
  CENX1 U2125 ( .A(n1588), .B(n1805), .Z(n1311) );
  CIVX2 U2126 ( .A(n1782), .Z(n1783) );
  CENX1 U2127 ( .A(n1831), .B(n1807), .Z(n1309) );
  CEOX1 U2128 ( .A(n329), .B(n147), .Z(product[3]) );
  CND2XL U2129 ( .A(n365), .B(n328), .Z(n147) );
  CNIVX1 U2130 ( .A(n830), .Z(n1778) );
  CEO3X1 U2131 ( .A(n403), .B(n1714), .C(n1715), .Z(n374) );
  CEN3X1 U2132 ( .A(n909), .B(n849), .C(n819), .Z(n1714) );
  CEN3X2 U2133 ( .A(n861), .B(n891), .C(n1059), .Z(n1715) );
  CEOX1 U2134 ( .A(n803), .B(n825), .Z(n382) );
  COR2X1 U2135 ( .A(n1716), .B(n1717), .Z(n966) );
  CAN2X1 U2136 ( .A(n383), .B(n368), .Z(n1718) );
  CNR2X1 U2137 ( .A(n383), .B(n368), .Z(n150) );
  CENX1 U2138 ( .A(n1831), .B(n1393), .Z(n1296) );
  CENX1 U2139 ( .A(n1854), .B(n1393), .Z(n1171) );
  CENX1 U2140 ( .A(n1842), .B(n1391), .Z(n1238) );
  CENX1 U2141 ( .A(n1837), .B(n1391), .Z(n1265) );
  CENX1 U2142 ( .A(n1831), .B(n1388), .Z(n1291) );
  CENX1 U2143 ( .A(n1588), .B(n1391), .Z(n1294) );
  CENX1 U2144 ( .A(n1833), .B(b[25]), .Z(n1258) );
  CENX1 U2145 ( .A(n1833), .B(n1388), .Z(n1262) );
  CENX1 U2146 ( .A(n104), .B(a[28]), .Z(n110) );
  CENX1 U2147 ( .A(n1839), .B(n1388), .Z(n1235) );
  CENX1 U2148 ( .A(n1819), .B(b[25]), .Z(n1318) );
  CENX1 U2149 ( .A(n1824), .B(b[24]), .Z(n1319) );
  CENX1 U2150 ( .A(n1824), .B(n1386), .Z(n1320) );
  CENX1 U2151 ( .A(n1843), .B(n1393), .Z(n1240) );
  CIVX4 U2152 ( .A(a[0]), .Z(n6) );
  CENX1 U2153 ( .A(n1831), .B(b[26]), .Z(n1286) );
  CENX1 U2154 ( .A(n1588), .B(b[24]), .Z(n1288) );
  CENX1 U2155 ( .A(n1820), .B(n1389), .Z(n1323) );
  CIVX2 U2156 ( .A(n12), .Z(n1825) );
  CND2XL U2157 ( .A(n1713), .B(n333), .Z(n148) );
  CENX1 U2158 ( .A(n1831), .B(b[27]), .Z(n1285) );
  CNIVX4 U2159 ( .A(n116), .Z(n1876) );
  CEOXL U2160 ( .A(a[30]), .B(a[31]), .Z(n1410) );
  CNIVX2 U2161 ( .A(n1397), .Z(n1815) );
  CHA1XL U2162 ( .A(n807), .B(n869), .CO(n581), .S(n582) );
  CNIVX1 U2163 ( .A(n66), .Z(n1776) );
  CIVX1 U2164 ( .A(n1859), .Z(n1779) );
  CIVXL U2165 ( .A(n1861), .Z(n1859) );
  CNR2IXL U2166 ( .B(n1876), .A(n58), .Z(n928) );
  CENX1 U2167 ( .A(n1860), .B(n1814), .Z(n1157) );
  COND2XL U2168 ( .A(n1619), .B(n1303), .C(n1302), .D(n24), .Z(n1018) );
  COND2XL U2169 ( .A(n1620), .B(n1312), .C(n1311), .D(n24), .Z(n1027) );
  COND2XL U2170 ( .A(n1619), .B(n1310), .C(n1309), .D(n24), .Z(n1025) );
  COND2XL U2171 ( .A(n1619), .B(n1587), .C(n1313), .D(n24), .Z(n816) );
  CFA1XL U2172 ( .A(n903), .B(n1013), .CI(n987), .CO(n651), .S(n652) );
  CNR2X1 U2173 ( .A(n248), .B(n251), .Z(n246) );
  CND2XL U2174 ( .A(n1773), .B(n1770), .Z(n133) );
  CNR2X1 U2175 ( .A(n1726), .B(n1724), .Z(n242) );
  CND2X1 U2176 ( .A(n1723), .B(n1722), .Z(n249) );
  CIVX2 U2177 ( .A(n1838), .Z(n1835) );
  CIVX2 U2178 ( .A(n30), .Z(n1838) );
  CENX1 U2179 ( .A(n1834), .B(n1809), .Z(n1278) );
  CFA1XL U2180 ( .A(n918), .B(n984), .CI(n938), .CO(n595), .S(n596) );
  COND2X1 U2181 ( .A(n107), .B(n1100), .C(n105), .D(n1099), .Z(n826) );
  CIVX1 U2182 ( .A(n1856), .Z(n1854) );
  CIVX1 U2183 ( .A(n1856), .Z(n1853) );
  CND2IXL U2184 ( .B(n1876), .A(n1852), .Z(n1188) );
  CFA1X1 U2185 ( .A(n1563), .B(n537), .CI(n956), .CO(n505), .S(n506) );
  COND2XL U2186 ( .A(n77), .B(n1861), .C(n1169), .D(n1639), .Z(n810) );
  CND2XL U2187 ( .A(net180512), .B(net179703), .Z(n127) );
  CIVX2 U2188 ( .A(n93), .Z(n1782) );
  COND2X1 U2189 ( .A(n1572), .B(n1128), .C(n1127), .D(n1651), .Z(n851) );
  CND2IXL U2190 ( .B(n1876), .A(n1583), .Z(n1209) );
  CENX1 U2191 ( .A(n1868), .B(n1810), .Z(n1130) );
  CENX1 U2192 ( .A(n1868), .B(n1809), .Z(n1131) );
  CND2IXL U2193 ( .B(n1876), .A(n1868), .Z(n1137) );
  COND2XL U2194 ( .A(n1620), .B(n1298), .C(n1297), .D(n24), .Z(n1013) );
  COND2XL U2195 ( .A(n27), .B(n1299), .C(n1298), .D(n24), .Z(n1014) );
  CNR2IXL U2196 ( .B(n1876), .A(n24), .Z(n1028) );
  COND2XL U2197 ( .A(n1620), .B(n1309), .C(n1308), .D(n24), .Z(n1024) );
  COND2XL U2198 ( .A(n1620), .B(n1305), .C(n1304), .D(n24), .Z(n1020) );
  COND2XL U2199 ( .A(n27), .B(n1289), .C(n1288), .D(n24), .Z(n1004) );
  COND2XL U2200 ( .A(n1619), .B(n1286), .C(n1285), .D(n24), .Z(n1001) );
  COND2X1 U2201 ( .A(n1620), .B(n1294), .C(n1293), .D(n24), .Z(n1009) );
  CND2XL U2202 ( .A(n902), .B(n1012), .Z(n1785) );
  CND2XL U2203 ( .A(n1016), .B(n990), .Z(n1791) );
  CFA1XL U2204 ( .A(n998), .B(n1024), .CI(n974), .CO(n783), .S(n784) );
  CIVXL U2205 ( .A(n1783), .Z(n1784) );
  CND2XL U2206 ( .A(n902), .B(n1070), .Z(n1786) );
  CND2XL U2207 ( .A(n1012), .B(n1070), .Z(n1787) );
  CND3X1 U2208 ( .A(n1785), .B(n1786), .C(n1787), .Z(n637) );
  CIVXL U2209 ( .A(n1583), .Z(n1788) );
  CFA1X1 U2210 ( .A(n850), .B(n862), .CI(n1002), .CO(n405), .S(n406) );
  COND2X1 U2211 ( .A(n1572), .B(n1127), .C(n1126), .D(n1650), .Z(n850) );
  COND2XL U2212 ( .A(n18), .B(n1324), .C(n1323), .D(n1574), .Z(n1038) );
  CND2XL U2213 ( .A(n966), .B(n1016), .Z(n1789) );
  CND2XL U2214 ( .A(n966), .B(n990), .Z(n1790) );
  CIVX2 U2215 ( .A(a[4]), .Z(n1793) );
  CND2X1 U2216 ( .A(n1821), .B(n1793), .Z(n1794) );
  CIVXL U2217 ( .A(n1835), .Z(n1797) );
  CND2IXL U2218 ( .B(n1876), .A(n1836), .Z(n1284) );
  CENX1 U2219 ( .A(n1834), .B(n1807), .Z(n1280) );
  CND2IXL U2220 ( .B(n1876), .A(n1849), .Z(n1232) );
  COND2XL U2221 ( .A(n61), .B(n1190), .C(n1189), .D(n58), .Z(n909) );
  COND2XL U2222 ( .A(n61), .B(n1191), .C(n1190), .D(n58), .Z(n910) );
  COND2XL U2223 ( .A(n61), .B(n1204), .C(n1203), .D(n58), .Z(n923) );
  COND2XL U2224 ( .A(n61), .B(n1193), .C(n1192), .D(n58), .Z(n912) );
  COND2XL U2225 ( .A(n61), .B(n1199), .C(n1198), .D(n58), .Z(n918) );
  COND2XL U2226 ( .A(n61), .B(n1198), .C(n1197), .D(n58), .Z(n917) );
  CIVX1 U2227 ( .A(n39), .Z(n1847) );
  CEOXL U2228 ( .A(n313), .B(n143), .Z(product[7]) );
  CNR2IXL U2229 ( .B(n1876), .A(n105), .Z(n830) );
  CANR1X2 U2230 ( .A(n1772), .B(n1753), .C(n269), .Z(n267) );
  CIVX2 U2231 ( .A(n1872), .Z(n1870) );
  CND2IXL U2232 ( .B(n1876), .A(n104), .Z(n1104) );
  CIVX1 U2233 ( .A(n1587), .Z(n1828) );
  CFA1X1 U2234 ( .A(n854), .B(n1006), .CI(n880), .CO(n511), .S(n512) );
  COND2X1 U2235 ( .A(n91), .B(n1131), .C(n1130), .D(n1651), .Z(n854) );
  COND2XL U2236 ( .A(n1654), .B(n1245), .C(n1244), .D(n1575), .Z(n962) );
  CIVX2 U2237 ( .A(n39), .Z(n1846) );
  COND2XL U2238 ( .A(n1559), .B(n1211), .C(n1210), .D(n1560), .Z(n929) );
  COND2XL U2239 ( .A(n1559), .B(n1212), .C(n1211), .D(n1557), .Z(n930) );
  COND2XL U2240 ( .A(n1559), .B(n1218), .C(n1217), .D(n1557), .Z(n936) );
  COND2XL U2241 ( .A(n1559), .B(n1227), .C(n1226), .D(n50), .Z(n945) );
  COND2XL U2242 ( .A(n1559), .B(n1225), .C(n1224), .D(n50), .Z(n943) );
  COND2XL U2243 ( .A(n1558), .B(n1221), .C(n1220), .D(n1560), .Z(n939) );
  COND2XL U2244 ( .A(n1559), .B(n1219), .C(n1218), .D(n50), .Z(n937) );
  COND2XL U2245 ( .A(n53), .B(n1231), .C(n1230), .D(n50), .Z(n949) );
  COND2XL U2246 ( .A(n1559), .B(n1220), .C(n1219), .D(n50), .Z(n938) );
  COND2XL U2247 ( .A(n1559), .B(n1222), .C(n1221), .D(n50), .Z(n940) );
  COND2XL U2248 ( .A(n1558), .B(n1224), .C(n1223), .D(n50), .Z(n942) );
  COND2XL U2249 ( .A(n1558), .B(n1216), .C(n1215), .D(n50), .Z(n934) );
  COND2XL U2250 ( .A(n1558), .B(n1229), .C(n1228), .D(n50), .Z(n947) );
  COND2XL U2251 ( .A(n1558), .B(n1223), .C(n1222), .D(n50), .Z(n941) );
  CNR2IX1 U2252 ( .B(n1876), .A(n110), .Z(n824) );
  COND2XL U2253 ( .A(n112), .B(n1436), .C(n110), .D(n1097), .Z(n804) );
  CND2X1 U2254 ( .A(n516), .B(n539), .Z(n193) );
  CND2XL U2255 ( .A(n1732), .B(n1731), .Z(n1800) );
  CND2X1 U2256 ( .A(n1732), .B(n1730), .Z(n1801) );
  CND2XL U2257 ( .A(n1731), .B(n1730), .Z(n1802) );
  CND3XL U2258 ( .A(n1800), .B(n1801), .C(n1802), .Z(n539) );
  CNR2X1 U2259 ( .A(n516), .B(n539), .Z(n192) );
  COAN1X1 U2260 ( .A(n243), .B(n1683), .C(n238), .Z(n234) );
  CENX1 U2261 ( .A(n1863), .B(n1806), .Z(n1149) );
  COND2XL U2262 ( .A(n36), .B(n1282), .C(n1281), .D(n1796), .Z(n998) );
  CNR2IXL U2263 ( .B(n1876), .A(n1796), .Z(n1000) );
  COND2XL U2264 ( .A(n1570), .B(n1267), .C(n1266), .D(n1796), .Z(n983) );
  COND2XL U2265 ( .A(n1570), .B(n1271), .C(n1270), .D(n1796), .Z(n987) );
  CND2X1 U2266 ( .A(n440), .B(n465), .Z(n172) );
  COND2XL U2267 ( .A(n1559), .B(n1595), .C(n1232), .D(n50), .Z(n813) );
  COND2XL U2268 ( .A(n1571), .B(n1259), .C(n1258), .D(n1796), .Z(n975) );
  COND2XL U2269 ( .A(n1570), .B(n1261), .C(n1260), .D(n1796), .Z(n977) );
  COND2XL U2270 ( .A(n1570), .B(n1281), .C(n1280), .D(n1796), .Z(n997) );
  COND2XL U2271 ( .A(n1571), .B(n1260), .C(n1259), .D(n1796), .Z(n976) );
  COND2XL U2272 ( .A(n1570), .B(n1279), .C(n1278), .D(n1796), .Z(n995) );
  COND2XL U2273 ( .A(n1571), .B(n1597), .C(n1284), .D(n1796), .Z(n815) );
  COND2XL U2274 ( .A(n1571), .B(n1283), .C(n1282), .D(n1796), .Z(n999) );
  COND2XL U2275 ( .A(n18), .B(n1568), .C(n1344), .D(n1573), .Z(n817) );
  CENX1 U2276 ( .A(n1819), .B(n1817), .Z(n1329) );
  CENX1 U2277 ( .A(n1833), .B(n1389), .Z(n1263) );
  CIVX1 U2278 ( .A(n1825), .Z(n1819) );
  CIVX1 U2279 ( .A(n1825), .Z(n1820) );
  CND2IXL U2280 ( .B(n1876), .A(n1823), .Z(n1344) );
  CENX1 U2281 ( .A(n1839), .B(n1390), .Z(n1237) );
  CENX1 U2282 ( .A(n1839), .B(n1389), .Z(n1236) );
  CIVX2 U2283 ( .A(n1845), .Z(n1839) );
  CANR1X2 U2284 ( .A(n261), .B(n1773), .C(n254), .Z(n252) );
  CIVX1 U2285 ( .A(n1587), .Z(n1826) );
  CENX1 U2286 ( .A(n1780), .B(n1811), .Z(n1161) );
  COND2X1 U2287 ( .A(n1572), .B(n1130), .C(n1129), .D(n1651), .Z(n853) );
  CANR1X2 U2288 ( .A(n246), .B(n1602), .C(n247), .Z(n245) );
  COND2XL U2289 ( .A(n1572), .B(n1126), .C(n1125), .D(n1650), .Z(n849) );
  CNR2IXL U2290 ( .B(n1876), .A(n1651), .Z(n860) );
  CND2IXL U2291 ( .B(n1876), .A(n1862), .Z(n1152) );
  CND2X4 U2292 ( .A(n1424), .B(n1590), .Z(n18) );
  CIVXL U2293 ( .A(n1825), .Z(n1822) );
  CIVXL U2294 ( .A(n1825), .Z(n1823) );
  CIVXL U2295 ( .A(n1587), .Z(n1827) );
  CIVXL U2296 ( .A(n1587), .Z(n1830) );
  CIVXL U2297 ( .A(n39), .Z(n1845) );
  CIVX2 U2298 ( .A(n327), .Z(n365) );
  CIVX2 U2299 ( .A(n319), .Z(n363) );
  CIVX2 U2300 ( .A(n248), .Z(n350) );
  CIVX2 U2301 ( .A(n333), .Z(n331) );
  CIVX2 U2302 ( .A(n325), .Z(n323) );
  CIVX2 U2303 ( .A(n317), .Z(n315) );
  CIVX2 U2304 ( .A(n309), .Z(n307) );
  CIVX2 U2305 ( .A(n303), .Z(n301) );
  CIVX2 U2306 ( .A(n1764), .Z(n279) );
  CIVX2 U2307 ( .A(n280), .Z(n355) );
  CIVX2 U2308 ( .A(n1769), .Z(n352) );
  CIVX2 U2309 ( .A(n242), .Z(n349) );
  CIVX2 U2310 ( .A(n156), .Z(n154) );
  CIVX2 U2311 ( .A(n109), .Z(n1436) );
endmodule


module calc_DW02_mult_2_stage_2 ( A, B, TC, CLK, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC, CLK;
  wire   n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, \A_extended[32] ,
         \B_extended[32] ;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33;
  assign \A_extended[32]  = A[31];
  assign \B_extended[32]  = B[31];

  calc_DW_mult_tc_25 mult_96 ( .a({\A_extended[32] , \A_extended[32] , A[30:2], 
        1'b0, A[0]}), .b({\B_extended[32] , \B_extended[32] , B[30:0]}), 
        .product({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, PRODUCT[31:10], 
        n16, n17, n18, n19, n20, n21, n22, n23, n24, n25}), 
        .i_retiming_group_0_clk(CLK) );
  CFD1QX1 clk_r_REG282_S1 ( .D(n16), .CP(CLK), .Q(PRODUCT[9]) );
  CFD1QX1 clk_r_REG344_S1 ( .D(n17), .CP(CLK), .Q(PRODUCT[8]) );
  CFD1QX1 clk_r_REG346_S1 ( .D(n19), .CP(CLK), .Q(PRODUCT[6]) );
  CFD1QX1 clk_r_REG348_S1 ( .D(n21), .CP(CLK), .Q(PRODUCT[4]) );
  CFD1QX1 clk_r_REG349_S1 ( .D(n22), .CP(CLK), .Q(PRODUCT[3]) );
  CFD1QX1 clk_r_REG352_S1 ( .D(n25), .CP(CLK), .Q(PRODUCT[0]) );
  CFD1QX4 clk_r_REG351_S1 ( .D(n24), .CP(CLK), .Q(PRODUCT[1]) );
  CFD1QX4 clk_r_REG347_S1 ( .D(n20), .CP(CLK), .Q(PRODUCT[5]) );
  CFD1QX4 clk_r_REG350_S1 ( .D(n23), .CP(CLK), .Q(PRODUCT[2]) );
  CFD1QX2 clk_r_REG345_S1 ( .D(n18), .CP(CLK), .Q(PRODUCT[7]) );
endmodule


module calc_DW_mult_tc_14 ( a, b, product, i_retiming_group_1_clk );
  input [32:0] a;
  input [32:0] b;
  output [65:0] product;
  input i_retiming_group_1_clk;
  wire   n6, n12, n15, n18, n21, n24, n27, n30, n36, n39, n42, n44, n48, n50,
         n53, n55, n58, n61, n63, n66, n69, n71, n74, n77, n79, n82, n84, n86,
         n89, n91, n93, n95, n97, n99, n100, n102, n104, n105, n107, n109,
         n110, n112, n113, n114, n115, n116, n121, n122, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n151,
         n152, n158, n160, n161, n163, n165, n166, n167, n168, n169, n170,
         n171, n172, n174, n175, n176, n179, n180, n181, n182, n184, n187,
         n188, n189, n191, n192, n193, n194, n195, n196, n197, n199, n201,
         n203, n204, n205, n206, n210, n212, n213, n214, n215, n216, n217,
         n221, n223, n224, n225, n226, n228, n231, n232, n233, n234, n236,
         n238, n239, n241, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n254, n256, n257, n258, n259, n261, n264, n265, n266,
         n267, n269, n271, n272, n273, n274, n275, n276, n277, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n296, n298, n299, n301, n303, n304, n305, n307,
         n309, n310, n311, n312, n313, n315, n317, n318, n319, n320, n321,
         n323, n325, n326, n327, n328, n329, n331, n333, n335, n340, n341,
         n342, n343, n347, n350, n352, n354, n355, n356, n357, n365, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1420,
         n1421, n1422, n1423, n1424, n1435, n1436, n1437, n1901, n1900, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899;
  assign n12 = a[3];
  assign n21 = a[5];
  assign n30 = a[7];
  assign n39 = a[9];
  assign n48 = a[11];
  assign n55 = a[13];
  assign n63 = a[15];
  assign n71 = a[17];
  assign n79 = a[19];
  assign n86 = a[21];
  assign n93 = a[23];
  assign n99 = a[25];
  assign n104 = a[27];
  assign n109 = a[29];
  assign n113 = a[32];
  assign n116 = b[0];
  assign n1386 = b[23];
  assign n1387 = b[22];
  assign n1388 = b[21];
  assign n1389 = b[20];
  assign n1390 = b[19];
  assign n1391 = b[18];
  assign n1392 = b[17];
  assign n1393 = b[16];
  assign n1394 = b[15];
  assign n1395 = b[14];
  assign n1396 = b[13];
  assign n1397 = b[12];
  assign n1398 = b[11];
  assign n1399 = b[10];
  assign n1400 = b[9];
  assign n1401 = b[8];
  assign n1402 = b[7];
  assign n1403 = b[6];
  assign n1404 = b[5];
  assign n1405 = b[4];
  assign n1406 = b[3];
  assign n1407 = b[2];
  assign n1408 = b[1];
  assign n1823 = i_retiming_group_1_clk;

  CEO3X2 U375 ( .A(n387), .B(n369), .C(n385), .Z(n368) );
  CEO3X2 U376 ( .A(n389), .B(n371), .C(n370), .Z(n369) );
  CEO3X2 U377 ( .A(n373), .B(n391), .C(n372), .Z(n370) );
  CEO3X2 U378 ( .A(n374), .B(n375), .C(n393), .Z(n371) );
  CEO3X2 U379 ( .A(n1815), .B(n397), .C(n395), .Z(n372) );
  CEO3X2 U380 ( .A(n1813), .B(n1814), .C(n1792), .Z(n373) );
  CEO3X2 U381 ( .A(n1810), .B(n1786), .C(n1812), .Z(n374) );
  CEO3X2 U382 ( .A(n1811), .B(n1788), .C(n1790), .Z(n375) );
  CEO3X2 U383 ( .A(n409), .B(n382), .C(n407), .Z(n376) );
  CEO3X2 U385 ( .A(n891), .B(n975), .C(n1029), .Z(n378) );
  CEO3X2 U387 ( .A(n803), .B(n849), .C(n861), .Z(n380) );
  CEO3X2 U388 ( .A(n821), .B(n819), .C(n839), .Z(n381) );
  CFA1X1 U390 ( .A(n388), .B(n386), .CI(n413), .CO(n383), .S(n384) );
  CFA1X1 U391 ( .A(n417), .B(n415), .CI(n390), .CO(n385), .S(n386) );
  CFA1X1 U392 ( .A(n394), .B(n392), .CI(n419), .CO(n387), .S(n388) );
  CFA1X1 U393 ( .A(n398), .B(n396), .CI(n421), .CO(n389), .S(n390) );
  CFA1X1 U394 ( .A(n425), .B(n423), .CI(n1791), .CO(n391), .S(n392) );
  CFA1X1 U395 ( .A(n1785), .B(n1789), .CI(n1787), .CO(n393), .S(n394) );
  CFA1X1 U396 ( .A(n1778), .B(n1782), .CI(n1784), .CO(n395), .S(n396) );
  CFA1X1 U397 ( .A(n1776), .B(n1780), .CI(n1783), .CO(n397), .S(n398) );
  CFA1X1 U398 ( .A(n952), .B(n435), .CI(n437), .CO(n399), .S(n400) );
  CFA1X1 U399 ( .A(n910), .B(n1060), .CI(n976), .CO(n401), .S(n402) );
  CFA1X1 U401 ( .A(n862), .B(n1002), .CI(n892), .CO(n405), .S(n406) );
  CFA1X1 U402 ( .A(n832), .B(n850), .CI(n840), .CO(n407), .S(n408) );
  CFA1X1 U403 ( .A(n820), .B(n822), .CI(n826), .CO(n409), .S(n410) );
  CFA1X1 U404 ( .A(n416), .B(n414), .CI(n441), .CO(n411), .S(n412) );
  CFA1X1 U405 ( .A(n420), .B(n443), .CI(n418), .CO(n413), .S(n414) );
  CFA1X1 U406 ( .A(n422), .B(n445), .CI(n447), .CO(n415), .S(n416) );
  CFA1X1 U407 ( .A(n426), .B(n424), .CI(n449), .CO(n417), .S(n418) );
  CFA1X1 U408 ( .A(n1781), .B(n451), .CI(n453), .CO(n419), .S(n420) );
  CFA1X1 U409 ( .A(n1775), .B(n1779), .CI(n1777), .CO(n421), .S(n422) );
  CFA1X1 U410 ( .A(n1773), .B(n1774), .CI(n1771), .CO(n423), .S(n424) );
  CFA1X1 U411 ( .A(n1765), .B(n1769), .CI(n1767), .CO(n425), .S(n426) );
  CFA1X1 U412 ( .A(n953), .B(n438), .CI(n1061), .CO(n427), .S(n428) );
  CFA1X1 U413 ( .A(n893), .B(n1003), .CI(n977), .CO(n429), .S(n430) );
  CFA1X1 U414 ( .A(n877), .B(n1031), .CI(n931), .CO(n431), .S(n432) );
  CFA1X1 U415 ( .A(n851), .B(n911), .CI(n863), .CO(n433), .S(n434) );
  CFA1X1 U416 ( .A(n804), .B(n841), .CI(n823), .CO(n435), .S(n436) );
  CHA1X1 U417 ( .A(n827), .B(n833), .CO(n437), .S(n438) );
  CFA1X1 U419 ( .A(n448), .B(n469), .CI(n446), .CO(n441), .S(n442) );
  CFA1X1 U420 ( .A(n450), .B(n471), .CI(n473), .CO(n443), .S(n444) );
  CFA1X1 U421 ( .A(n475), .B(n452), .CI(n454), .CO(n445), .S(n446) );
  CFA1X1 U422 ( .A(n1772), .B(n477), .CI(n1763), .CO(n447), .S(n448) );
  CFA1X1 U423 ( .A(n1766), .B(n1770), .CI(n1768), .CO(n449), .S(n450) );
  CFA1X1 U424 ( .A(n1757), .B(n1761), .CI(n1759), .CO(n451), .S(n452) );
  CFA1X1 U425 ( .A(n1809), .B(n1764), .CI(n1755), .CO(n453), .S(n454) );
  CFA1X1 U426 ( .A(n912), .B(n1062), .CI(n954), .CO(n455), .S(n456) );
  CFA1X1 U427 ( .A(n894), .B(n1032), .CI(n978), .CO(n457), .S(n458) );
  CFA1X1 U428 ( .A(n878), .B(n1004), .CI(n932), .CO(n459), .S(n460) );
  CFA1X1 U429 ( .A(n842), .B(n864), .CI(n852), .CO(n461), .S(n462) );
  CFA1X1 U430 ( .A(n824), .B(n834), .CI(n828), .CO(n463), .S(n464) );
  CFA1X1 U431 ( .A(n470), .B(n468), .CI(n493), .CO(n465), .S(n466) );
  CFA1X1 U432 ( .A(n497), .B(n495), .CI(n472), .CO(n467), .S(n468) );
  CFA1X1 U433 ( .A(n499), .B(n474), .CI(n476), .CO(n469), .S(n470) );
  CFA1X1 U434 ( .A(n503), .B(n478), .CI(n501), .CO(n471), .S(n472) );
  CFA1X1 U435 ( .A(n1758), .B(n1762), .CI(n1760), .CO(n473), .S(n474) );
  CFA1X1 U436 ( .A(n1753), .B(n1756), .CI(n1754), .CO(n475), .S(n476) );
  CFA1X1 U437 ( .A(n1747), .B(n1751), .CI(n1749), .CO(n477), .S(n478) );
  CFA1X1 U438 ( .A(n513), .B(n955), .CI(n490), .CO(n479), .S(n480) );
  CFA1X1 U439 ( .A(n913), .B(n979), .CI(n1063), .CO(n481), .S(n482) );
  CFA1X1 U441 ( .A(n865), .B(n1033), .CI(n895), .CO(n485), .S(n486) );
  CFA1X1 U442 ( .A(n829), .B(n853), .CI(n843), .CO(n487), .S(n488) );
  CHA1X1 U443 ( .A(n805), .B(n835), .CO(n489), .S(n490) );
  CFA1X1 U444 ( .A(n496), .B(n494), .CI(n517), .CO(n491), .S(n492) );
  CFA1X1 U445 ( .A(n521), .B(n519), .CI(n498), .CO(n493), .S(n494) );
  CFA1X1 U446 ( .A(n523), .B(n500), .CI(n502), .CO(n495), .S(n496) );
  CFA1X1 U447 ( .A(n527), .B(n504), .CI(n525), .CO(n497), .S(n498) );
  CFA1X1 U448 ( .A(n1748), .B(n1752), .CI(n1750), .CO(n499), .S(n500) );
  CFA1X1 U449 ( .A(n1742), .B(n1746), .CI(n1745), .CO(n501), .S(n502) );
  CFA1X1 U450 ( .A(n1738), .B(n1744), .CI(n1740), .CO(n503), .S(n504) );
  CFA1X1 U451 ( .A(n956), .B(n537), .CI(n1064), .CO(n505), .S(n506) );
  CFA1X1 U452 ( .A(n896), .B(n1006), .CI(n980), .CO(n507), .S(n508) );
  CFA1X1 U453 ( .A(n880), .B(n1034), .CI(n934), .CO(n509), .S(n510) );
  CFA1X1 U455 ( .A(n830), .B(n844), .CI(n836), .CO(n513), .S(n514) );
  CFA1X1 U456 ( .A(n520), .B(n518), .CI(n541), .CO(n515), .S(n516) );
  CFA1X1 U457 ( .A(n545), .B(n543), .CI(n522), .CO(n517), .S(n518) );
  CFA1X1 U458 ( .A(n547), .B(n524), .CI(n526), .CO(n519), .S(n520) );
  CFA1X1 U459 ( .A(n551), .B(n528), .CI(n549), .CO(n521), .S(n522) );
  CFA1X1 U460 ( .A(n1739), .B(n1743), .CI(n1741), .CO(n523), .S(n524) );
  CFA1X1 U461 ( .A(n1734), .B(n1737), .CI(n1736), .CO(n525), .S(n526) );
  CFA1X1 U462 ( .A(n1808), .B(n1732), .CI(n1730), .CO(n527), .S(n528) );
  CFA1X1 U463 ( .A(n915), .B(n1065), .CI(n957), .CO(n529), .S(n530) );
  CFA1X1 U465 ( .A(n881), .B(n1035), .CI(n935), .CO(n533), .S(n534) );
  CFA1X1 U466 ( .A(n845), .B(n867), .CI(n855), .CO(n535), .S(n536) );
  CHA1X1 U467 ( .A(n806), .B(n837), .CO(n537), .S(n538) );
  CFA1X1 U468 ( .A(n544), .B(n542), .CI(n563), .CO(n539), .S(n540) );
  CFA1X1 U470 ( .A(n569), .B(n548), .CI(n550), .CO(n543), .S(n544) );
  CFA1X1 U472 ( .A(n1731), .B(n1728), .CI(n1733), .CO(n547), .S(n548) );
  CFA1X1 U473 ( .A(n1724), .B(n1729), .CI(n1726), .CO(n549), .S(n550) );
  CFA1X1 U475 ( .A(n916), .B(n1066), .CI(n982), .CO(n553), .S(n554) );
  CFA1X1 U476 ( .A(n882), .B(n1036), .CI(n936), .CO(n555), .S(n556) );
  CFA1X1 U477 ( .A(n868), .B(n1008), .CI(n898), .CO(n557), .S(n558) );
  CFA1X1 U478 ( .A(n838), .B(n856), .CI(n846), .CO(n559), .S(n560) );
  CFA1X1 U482 ( .A(n1725), .B(n593), .CI(n1727), .CO(n567), .S(n568) );
  CFA1X1 U483 ( .A(n1718), .B(n1723), .CI(n1721), .CO(n569), .S(n570) );
  CFA1X1 U484 ( .A(n1714), .B(n1720), .CI(n1716), .CO(n571), .S(n572) );
  CFA1X1 U485 ( .A(n937), .B(n582), .CI(n959), .CO(n573), .S(n574) );
  CFA1X1 U486 ( .A(n917), .B(n1009), .CI(n1067), .CO(n575), .S(n576) );
  CHA1X1 U489 ( .A(n807), .B(n857), .CO(n581), .S(n582) );
  CFA1X1 U490 ( .A(n588), .B(n586), .CI(n605), .CO(n583), .S(n584) );
  CFA1X1 U491 ( .A(n592), .B(n607), .CI(n590), .CO(n585), .S(n586) );
  CFA1X1 U492 ( .A(n611), .B(n609), .CI(n594), .CO(n587), .S(n588) );
  CFA1X1 U494 ( .A(n1712), .B(n1715), .CI(n1713), .CO(n591), .S(n592) );
  CFA1X1 U495 ( .A(n1806), .B(n1710), .CI(n1708), .CO(n593), .S(n594) );
  CFA1X1 U496 ( .A(n918), .B(n1068), .CI(n960), .CO(n595), .S(n596) );
  CFA1X1 U497 ( .A(n900), .B(n1038), .CI(n984), .CO(n597), .S(n598) );
  CFA1X1 U498 ( .A(n884), .B(n1010), .CI(n938), .CO(n599), .S(n600) );
  CFA1X1 U500 ( .A(n608), .B(n606), .CI(n625), .CO(n603), .S(n604) );
  CFA1X1 U501 ( .A(n612), .B(n627), .CI(n610), .CO(n605), .S(n606) );
  CFA1X1 U502 ( .A(n631), .B(n629), .CI(n614), .CO(n607), .S(n608) );
  CFA1X1 U503 ( .A(n1706), .B(n1711), .CI(n1709), .CO(n609), .S(n610) );
  CFA1X1 U504 ( .A(n1702), .B(n1707), .CI(n1704), .CO(n611), .S(n612) );
  CFA1X1 U506 ( .A(n939), .B(n1039), .CI(n1069), .CO(n615), .S(n616) );
  CFA1X1 U507 ( .A(n901), .B(n1011), .CI(n985), .CO(n617), .S(n618) );
  CFA1X1 U508 ( .A(n859), .B(n919), .CI(n885), .CO(n619), .S(n620) );
  CHA1X1 U509 ( .A(n808), .B(n871), .CO(n621), .S(n622) );
  CFA1X1 U510 ( .A(n628), .B(n626), .CI(n643), .CO(n623), .S(n624) );
  CFA1X1 U511 ( .A(n632), .B(n645), .CI(n630), .CO(n625), .S(n626) );
  CFA1X1 U512 ( .A(n1705), .B(n647), .CI(n649), .CO(n627), .S(n628) );
  CFA1X1 U513 ( .A(n1699), .B(n1703), .CI(n1701), .CO(n629), .S(n630) );
  CFA1X1 U514 ( .A(n1694), .B(n1696), .CI(n1698), .CO(n631), .S(n632) );
  CFA1X1 U515 ( .A(n940), .B(n657), .CI(n962), .CO(n633), .S(n634) );
  CFA1X1 U516 ( .A(n920), .B(n1012), .CI(n1070), .CO(n635), .S(n636) );
  CFA1X1 U517 ( .A(n902), .B(n1040), .CI(n986), .CO(n637), .S(n638) );
  CFA1X1 U519 ( .A(n646), .B(n644), .CI(n661), .CO(n641), .S(n642) );
  CFA1X1 U520 ( .A(n650), .B(n663), .CI(n648), .CO(n643), .S(n644) );
  CFA1X1 U521 ( .A(n1697), .B(n665), .CI(n667), .CO(n645), .S(n646) );
  CFA1X1 U522 ( .A(n1690), .B(n1695), .CI(n1693), .CO(n647), .S(n648) );
  CFA1X1 U523 ( .A(n1804), .B(n1692), .CI(n1688), .CO(n649), .S(n650) );
  CFA1X1 U524 ( .A(n941), .B(n987), .CI(n963), .CO(n651), .S(n652) );
  CFA1X1 U525 ( .A(n921), .B(n1071), .CI(n1041), .CO(n653), .S(n654) );
  CFA1X1 U526 ( .A(n873), .B(n1013), .CI(n887), .CO(n655), .S(n656) );
  CHA1X1 U527 ( .A(n809), .B(n903), .CO(n657), .S(n658) );
  CFA1X1 U528 ( .A(n664), .B(n662), .CI(n677), .CO(n659), .S(n660) );
  CFA1X1 U529 ( .A(n668), .B(n679), .CI(n666), .CO(n661), .S(n662) );
  CFA1X1 U530 ( .A(n1691), .B(n681), .CI(n683), .CO(n663), .S(n664) );
  CFA1X1 U531 ( .A(n1686), .B(n1689), .CI(n1687), .CO(n665), .S(n666) );
  CFA1X1 U532 ( .A(n1637), .B(n1684), .CI(n1803), .CO(n667), .S(n668) );
  CFA1X1 U533 ( .A(n942), .B(n1072), .CI(n988), .CO(n669), .S(n670) );
  CFA1X1 U535 ( .A(n874), .B(n904), .CI(n888), .CO(n673), .S(n674) );
  CFA1X1 U536 ( .A(n680), .B(n678), .CI(n693), .CO(n675), .S(n676) );
  CFA1X1 U537 ( .A(n684), .B(n695), .CI(n682), .CO(n677), .S(n678) );
  CFA1X1 U538 ( .A(n1683), .B(n697), .CI(n1685), .CO(n679), .S(n680) );
  CFA1X1 U539 ( .A(n1678), .B(n1682), .CI(n1680), .CO(n681), .S(n682) );
  CFA1X1 U540 ( .A(n1641), .B(n1802), .CI(n1633), .CO(n683), .S(n684) );
  CFA1X1 U542 ( .A(n889), .B(n1043), .CI(n943), .CO(n687), .S(n688) );
  CHA1X1 U543 ( .A(n810), .B(n965), .CO(n689), .S(n690) );
  CFA1X1 U544 ( .A(n696), .B(n694), .CI(n707), .CO(n691), .S(n692) );
  CFA1X1 U545 ( .A(n711), .B(n709), .CI(n698), .CO(n693), .S(n694) );
  CFA1X1 U546 ( .A(n1677), .B(n1681), .CI(n1679), .CO(n695), .S(n696) );
  CFA1X1 U547 ( .A(n1801), .B(n1674), .CI(n1676), .CO(n697), .S(n698) );
  CFA1X1 U548 ( .A(n966), .B(n1074), .CI(n990), .CO(n699), .S(n700) );
  CFA1X1 U549 ( .A(n944), .B(n1044), .CI(n1016), .CO(n701), .S(n702) );
  CFA1X1 U550 ( .A(n890), .B(n924), .CI(n906), .CO(n703), .S(n704) );
  CFA1X1 U551 ( .A(n710), .B(n708), .CI(n721), .CO(n705), .S(n706) );
  CFA1X1 U552 ( .A(n1672), .B(n712), .CI(n723), .CO(n707), .S(n708) );
  CFA1X1 U553 ( .A(n1670), .B(n1675), .CI(n1673), .CO(n709), .S(n710) );
  CFA1X1 U554 ( .A(n1640), .B(n1668), .CI(n1800), .CO(n711), .S(n712) );
  CFA1X1 U555 ( .A(n925), .B(n1075), .CI(n967), .CO(n713), .S(n714) );
  CFA1X1 U556 ( .A(n907), .B(n1017), .CI(n991), .CO(n715), .S(n716) );
  CHA1X1 U557 ( .A(n811), .B(n1045), .CO(n717), .S(n718) );
  CFA1X1 U558 ( .A(n724), .B(n722), .CI(n733), .CO(n719), .S(n720) );
  CFA1X1 U559 ( .A(n1669), .B(n735), .CI(n1671), .CO(n721), .S(n722) );
  CFA1X1 U560 ( .A(n1666), .B(n1667), .CI(n1664), .CO(n723), .S(n724) );
  CFA1X1 U561 ( .A(n992), .B(n741), .CI(n1076), .CO(n725), .S(n726) );
  CFA1X1 U564 ( .A(n736), .B(n734), .CI(n745), .CO(n731), .S(n732) );
  CFA1X1 U565 ( .A(n1663), .B(n747), .CI(n1665), .CO(n733), .S(n734) );
  CFA1X1 U566 ( .A(n1799), .B(n1662), .CI(n1660), .CO(n735), .S(n736) );
  CFA1X1 U567 ( .A(n947), .B(n993), .CI(n969), .CO(n737), .S(n738) );
  CFA1X1 U568 ( .A(n927), .B(n1019), .CI(n1077), .CO(n739), .S(n740) );
  CHA1X1 U569 ( .A(n812), .B(n1047), .CO(n741), .S(n742) );
  CFA1X1 U570 ( .A(n755), .B(n746), .CI(n748), .CO(n743), .S(n744) );
  CFA1X1 U571 ( .A(n1659), .B(n757), .CI(n1661), .CO(n745), .S(n746) );
  CFA1X1 U572 ( .A(n1632), .B(n1658), .CI(n1798), .CO(n747), .S(n748) );
  CFA1X1 U573 ( .A(n994), .B(n1048), .CI(n1020), .CO(n749), .S(n750) );
  CFA1X1 U575 ( .A(n758), .B(n756), .CI(n765), .CO(n753), .S(n754) );
  CFA1X1 U576 ( .A(n1654), .B(n1657), .CI(n1656), .CO(n755), .S(n756) );
  CFA1X1 U577 ( .A(n1636), .B(n1797), .CI(n1631), .CO(n757), .S(n758) );
  CFA1X1 U578 ( .A(n949), .B(n1021), .CI(n1079), .CO(n759), .S(n760) );
  CHA1X1 U579 ( .A(n813), .B(n1049), .CO(n761), .S(n762) );
  CFA1X1 U580 ( .A(n1655), .B(n766), .CI(n773), .CO(n763), .S(n764) );
  CFA1X1 U581 ( .A(n1796), .B(n1653), .CI(n1652), .CO(n765), .S(n766) );
  CFA1X1 U582 ( .A(n1080), .B(n1050), .CI(n1022), .CO(n767), .S(n768) );
  CFA1X1 U583 ( .A(n950), .B(n996), .CI(n972), .CO(n769), .S(n770) );
  CFA1X1 U584 ( .A(n1650), .B(n774), .CI(n1651), .CO(n771), .S(n772) );
  CFA1X1 U585 ( .A(n1635), .B(n1648), .CI(n1795), .CO(n773), .S(n774) );
  CFA1X1 U586 ( .A(n973), .B(n1023), .CI(n1081), .CO(n775), .S(n776) );
  CHA1X1 U587 ( .A(n814), .B(n1051), .CO(n777), .S(n778) );
  CFA1X1 U588 ( .A(n1646), .B(n1649), .CI(n1647), .CO(n779), .S(n780) );
  CFA1X1 U589 ( .A(n1052), .B(n789), .CI(n1024), .CO(n781), .S(n782) );
  CFA1X1 U590 ( .A(n974), .B(n1082), .CI(n998), .CO(n783), .S(n784) );
  CFA1X1 U591 ( .A(n1794), .B(n1645), .CI(n1644), .CO(n785), .S(n786) );
  CFA1X1 U592 ( .A(n999), .B(n1025), .CI(n1083), .CO(n787), .S(n788) );
  CHA1X1 U593 ( .A(n815), .B(n1053), .CO(n789), .S(n790) );
  CFA1X1 U594 ( .A(n1634), .B(n1643), .CI(n1793), .CO(n791), .S(n792) );
  CFA1X1 U595 ( .A(n1000), .B(n1054), .CI(n1084), .CO(n793), .S(n794) );
  CFA1X1 U596 ( .A(n1055), .B(n798), .CI(n1027), .CO(n795), .S(n796) );
  CHA1X1 U597 ( .A(n1085), .B(n816), .CO(n797), .S(n798) );
  CFA1X1 U598 ( .A(n1028), .B(n1056), .CI(n1086), .CO(n799), .S(n800) );
  CHA1X1 U599 ( .A(n1087), .B(n1057), .CO(n801), .S(n802) );
  COND2X1 U600 ( .A(n115), .B(n1435), .C(n114), .D(n1092), .Z(n803) );
  COND2X1 U601 ( .A(n1091), .B(n115), .C(n114), .D(n1090), .Z(n819) );
  COND2X1 U606 ( .A(n112), .B(n1436), .C(n110), .D(n1097), .Z(n804) );
  COND2X1 U607 ( .A(n112), .B(n1094), .C(n110), .D(n1093), .Z(n821) );
  COND2X1 U608 ( .A(n112), .B(n1095), .C(n110), .D(n1094), .Z(n822) );
  COND2X1 U609 ( .A(n1096), .B(n112), .C(n110), .D(n1095), .Z(n823) );
  COND2X1 U630 ( .A(n102), .B(n1897), .C(n100), .D(n1113), .Z(n806) );
  COND2X1 U631 ( .A(n102), .B(n1106), .C(n1105), .D(n100), .Z(n831) );
  COND2X1 U632 ( .A(n102), .B(n1107), .C(n1106), .D(n100), .Z(n832) );
  COND2X1 U637 ( .A(n1112), .B(n102), .C(n1111), .D(n100), .Z(n837) );
  CND2IX1 U647 ( .B(n1899), .A(n1896), .Z(n1113) );
  COND2X1 U648 ( .A(n97), .B(n1895), .C(n1124), .D(n95), .Z(n807) );
  COND2X1 U649 ( .A(n97), .B(n1115), .C(n1114), .D(n95), .Z(n839) );
  COND2X1 U650 ( .A(n97), .B(n1116), .C(n1115), .D(n95), .Z(n840) );
  COND2X1 U651 ( .A(n97), .B(n1117), .C(n1116), .D(n95), .Z(n841) );
  COND2X1 U652 ( .A(n97), .B(n1118), .C(n1117), .D(n95), .Z(n842) );
  CND2IX1 U669 ( .B(n1899), .A(n1894), .Z(n1124) );
  COND2X1 U671 ( .A(n91), .B(n1126), .C(n1125), .D(n89), .Z(n849) );
  COND2X1 U672 ( .A(n91), .B(n1127), .C(n1126), .D(n89), .Z(n850) );
  COND2X1 U673 ( .A(n91), .B(n1128), .C(n1127), .D(n89), .Z(n851) );
  COND2X1 U674 ( .A(n91), .B(n1129), .C(n1128), .D(n89), .Z(n852) );
  COND2X1 U676 ( .A(n91), .B(n1131), .C(n1130), .D(n89), .Z(n854) );
  COND2X1 U677 ( .A(n91), .B(n1132), .C(n1131), .D(n89), .Z(n855) );
  COND2X1 U681 ( .A(n91), .B(n1136), .C(n1135), .D(n89), .Z(n859) );
  COND2X1 U696 ( .A(n84), .B(n1889), .C(n1152), .D(n82), .Z(n809) );
  COND2X1 U697 ( .A(n84), .B(n1139), .C(n1138), .D(n82), .Z(n861) );
  COND2X1 U698 ( .A(n84), .B(n1140), .C(n1139), .D(n82), .Z(n862) );
  COND2X1 U699 ( .A(n84), .B(n1141), .C(n1140), .D(n82), .Z(n863) );
  COND2X1 U700 ( .A(n84), .B(n1142), .C(n1141), .D(n82), .Z(n864) );
  COND2X1 U702 ( .A(n84), .B(n1144), .C(n1143), .D(n82), .Z(n866) );
  COND2X1 U703 ( .A(n84), .B(n1145), .C(n1144), .D(n82), .Z(n867) );
  COND2X1 U704 ( .A(n84), .B(n1146), .C(n1145), .D(n82), .Z(n868) );
  CND2IX1 U725 ( .B(n1899), .A(n1886), .Z(n1152) );
  COND2X1 U726 ( .A(n77), .B(n1885), .C(n1169), .D(n74), .Z(n810) );
  COND2X1 U727 ( .A(n77), .B(n1154), .C(n1153), .D(n74), .Z(n875) );
  COND2X1 U729 ( .A(n77), .B(n1156), .C(n1155), .D(n74), .Z(n877) );
  COND2X1 U730 ( .A(n77), .B(n1157), .C(n1156), .D(n74), .Z(n878) );
  COND2X1 U731 ( .A(n77), .B(n1158), .C(n1157), .D(n74), .Z(n879) );
  COND2X1 U732 ( .A(n77), .B(n1159), .C(n1158), .D(n74), .Z(n880) );
  COND2X1 U733 ( .A(n77), .B(n1160), .C(n1159), .D(n74), .Z(n881) );
  COND2X1 U734 ( .A(n77), .B(n1161), .C(n1160), .D(n74), .Z(n882) );
  COND2X1 U737 ( .A(n77), .B(n1164), .C(n1163), .D(n74), .Z(n885) );
  COND2X1 U741 ( .A(n77), .B(n1168), .C(n1167), .D(n74), .Z(n889) );
  CND2IX1 U759 ( .B(n1899), .A(n1882), .Z(n1169) );
  COND2X1 U761 ( .A(n69), .B(n1171), .C(n1170), .D(n66), .Z(n891) );
  COND2X1 U762 ( .A(n69), .B(n1172), .C(n1171), .D(n66), .Z(n892) );
  COND2X1 U763 ( .A(n69), .B(n1173), .C(n1172), .D(n66), .Z(n893) );
  COND2X1 U764 ( .A(n69), .B(n1174), .C(n1173), .D(n66), .Z(n894) );
  COND2X1 U766 ( .A(n69), .B(n1176), .C(n1175), .D(n66), .Z(n896) );
  COND2X1 U767 ( .A(n69), .B(n1177), .C(n1176), .D(n66), .Z(n897) );
  COND2X1 U768 ( .A(n69), .B(n1178), .C(n1177), .D(n66), .Z(n898) );
  COND2X1 U769 ( .A(n69), .B(n1179), .C(n1178), .D(n66), .Z(n899) );
  COND2X1 U771 ( .A(n69), .B(n1181), .C(n1180), .D(n66), .Z(n901) );
  COND2X1 U773 ( .A(n69), .B(n1183), .C(n1182), .D(n66), .Z(n903) );
  COND2X1 U774 ( .A(n69), .B(n1184), .C(n1183), .D(n66), .Z(n904) );
  COND2X1 U775 ( .A(n69), .B(n1185), .C(n1184), .D(n66), .Z(n905) );
  COND2X1 U776 ( .A(n69), .B(n1186), .C(n1185), .D(n66), .Z(n906) );
  COND2X1 U777 ( .A(n69), .B(n1187), .C(n1186), .D(n66), .Z(n907) );
  CND2IX1 U797 ( .B(n1899), .A(n1878), .Z(n1188) );
  COND2X1 U798 ( .A(n61), .B(n1877), .C(n1209), .D(n58), .Z(n812) );
  COND2X1 U799 ( .A(n61), .B(n1190), .C(n1189), .D(n58), .Z(n909) );
  COND2X1 U800 ( .A(n61), .B(n1191), .C(n1190), .D(n58), .Z(n910) );
  COND2X1 U801 ( .A(n61), .B(n1192), .C(n1191), .D(n58), .Z(n911) );
  COND2X1 U802 ( .A(n61), .B(n1193), .C(n1192), .D(n58), .Z(n912) );
  COND2X1 U803 ( .A(n61), .B(n1194), .C(n1193), .D(n58), .Z(n913) );
  COND2X1 U805 ( .A(n61), .B(n1196), .C(n1195), .D(n58), .Z(n915) );
  COND2X1 U806 ( .A(n61), .B(n1197), .C(n1196), .D(n58), .Z(n916) );
  COND2X1 U807 ( .A(n61), .B(n1198), .C(n1197), .D(n58), .Z(n917) );
  COND2X1 U815 ( .A(n61), .B(n1206), .C(n1205), .D(n58), .Z(n925) );
  COND2X1 U817 ( .A(n61), .B(n1208), .C(n1207), .D(n58), .Z(n927) );
  CND2IX1 U839 ( .B(n1899), .A(n1876), .Z(n1209) );
  COND2X1 U840 ( .A(n53), .B(n1874), .C(n1232), .D(n50), .Z(n813) );
  COND2X1 U841 ( .A(n53), .B(n1211), .C(n1210), .D(n50), .Z(n929) );
  COND2X1 U843 ( .A(n53), .B(n1213), .C(n1212), .D(n50), .Z(n931) );
  COND2X1 U847 ( .A(n53), .B(n1217), .C(n1216), .D(n50), .Z(n935) );
  COND2X1 U848 ( .A(n53), .B(n1218), .C(n1217), .D(n50), .Z(n936) );
  COND2X1 U850 ( .A(n53), .B(n1220), .C(n1219), .D(n50), .Z(n938) );
  COND2X1 U851 ( .A(n53), .B(n1221), .C(n1220), .D(n50), .Z(n939) );
  COND2X1 U852 ( .A(n53), .B(n1222), .C(n1221), .D(n50), .Z(n940) );
  COND2X1 U853 ( .A(n53), .B(n1223), .C(n1222), .D(n50), .Z(n941) );
  COND2X1 U854 ( .A(n53), .B(n1224), .C(n1223), .D(n50), .Z(n942) );
  COND2X1 U855 ( .A(n53), .B(n1225), .C(n1224), .D(n50), .Z(n943) );
  COND2X1 U856 ( .A(n53), .B(n1226), .C(n1225), .D(n50), .Z(n944) );
  COND2X1 U857 ( .A(n53), .B(n1227), .C(n1226), .D(n50), .Z(n945) );
  COND2X1 U859 ( .A(n53), .B(n1229), .C(n1228), .D(n50), .Z(n947) );
  COND2X1 U861 ( .A(n53), .B(n1231), .C(n1230), .D(n50), .Z(n949) );
  CND2IX1 U885 ( .B(n1899), .A(n1873), .Z(n1232) );
  COND2X1 U886 ( .A(n44), .B(n1871), .C(n1257), .D(n1836), .Z(n814) );
  COND2X1 U887 ( .A(n44), .B(n1234), .C(n1233), .D(n1836), .Z(n951) );
  COND2X1 U889 ( .A(n44), .B(n1236), .C(n1235), .D(n1836), .Z(n953) );
  COND2X1 U890 ( .A(n44), .B(n1237), .C(n1236), .D(n1836), .Z(n954) );
  COND2X1 U891 ( .A(n44), .B(n1238), .C(n1237), .D(n1836), .Z(n955) );
  COND2X1 U892 ( .A(n44), .B(n1239), .C(n1238), .D(n1836), .Z(n956) );
  COND2X1 U893 ( .A(n44), .B(n1240), .C(n1239), .D(n1836), .Z(n957) );
  COND2X1 U895 ( .A(n44), .B(n1242), .C(n1241), .D(n1836), .Z(n959) );
  COND2X1 U896 ( .A(n44), .B(n1243), .C(n1242), .D(n1836), .Z(n960) );
  COND2X1 U898 ( .A(n44), .B(n1245), .C(n1244), .D(n1836), .Z(n962) );
  COND2X1 U899 ( .A(n44), .B(n1246), .C(n1245), .D(n1836), .Z(n963) );
  COND2X1 U901 ( .A(n44), .B(n1248), .C(n1247), .D(n1836), .Z(n965) );
  COND2X1 U902 ( .A(n44), .B(n1249), .C(n1248), .D(n1836), .Z(n966) );
  COND2X1 U903 ( .A(n44), .B(n1250), .C(n1249), .D(n1836), .Z(n967) );
  COND2X1 U904 ( .A(n44), .B(n1251), .C(n1250), .D(n1836), .Z(n968) );
  COND2X1 U905 ( .A(n44), .B(n1252), .C(n1251), .D(n1836), .Z(n969) );
  COND2X1 U906 ( .A(n44), .B(n1253), .C(n1252), .D(n1836), .Z(n970) );
  COND2X1 U908 ( .A(n44), .B(n1255), .C(n1254), .D(n1836), .Z(n972) );
  COND2X1 U909 ( .A(n44), .B(n1256), .C(n1255), .D(n1836), .Z(n973) );
  CND2IX1 U935 ( .B(n1899), .A(n1867), .Z(n1257) );
  COND2X1 U936 ( .A(n36), .B(n1865), .C(n1284), .D(n1606), .Z(n815) );
  COND2X1 U937 ( .A(n1259), .B(n36), .C(n1258), .D(n1606), .Z(n975) );
  COND2X1 U941 ( .A(n36), .B(n1263), .C(n1262), .D(n1606), .Z(n979) );
  COND2X1 U942 ( .A(n36), .B(n1264), .C(n1263), .D(n1606), .Z(n980) );
  COND2X1 U945 ( .A(n36), .B(n1267), .C(n1266), .D(n1606), .Z(n983) );
  COND2X1 U946 ( .A(n36), .B(n1268), .C(n1267), .D(n1606), .Z(n984) );
  COND2X1 U949 ( .A(n36), .B(n1271), .C(n1270), .D(n1606), .Z(n987) );
  COND2X1 U950 ( .A(n36), .B(n1272), .C(n1271), .D(n1606), .Z(n988) );
  COND2X1 U951 ( .A(n36), .B(n1273), .C(n1272), .D(n1606), .Z(n989) );
  COND2X1 U952 ( .A(n36), .B(n1274), .C(n1273), .D(n1606), .Z(n990) );
  COND2X1 U953 ( .A(n36), .B(n1275), .C(n1274), .D(n1606), .Z(n991) );
  COND2X1 U954 ( .A(n36), .B(n1276), .C(n1275), .D(n1606), .Z(n992) );
  COND2X1 U955 ( .A(n36), .B(n1277), .C(n1276), .D(n1606), .Z(n993) );
  COND2X1 U956 ( .A(n36), .B(n1278), .C(n1277), .D(n1606), .Z(n994) );
  COND2X1 U959 ( .A(n36), .B(n1281), .C(n1280), .D(n1606), .Z(n997) );
  COND2X1 U961 ( .A(n36), .B(n1283), .C(n1282), .D(n1606), .Z(n999) );
  CND2IX1 U989 ( .B(n1899), .A(n1861), .Z(n1284) );
  COND2X1 U990 ( .A(n27), .B(n1860), .C(n1313), .D(n24), .Z(n816) );
  COND2X1 U992 ( .A(n27), .B(n1287), .C(n24), .D(n1286), .Z(n1002) );
  COND2X1 U993 ( .A(n27), .B(n1288), .C(n24), .D(n1287), .Z(n1003) );
  COND2X1 U994 ( .A(n27), .B(n1289), .C(n24), .D(n1288), .Z(n1004) );
  COND2X1 U995 ( .A(n27), .B(n1290), .C(n24), .D(n1289), .Z(n1005) );
  COND2X1 U996 ( .A(n27), .B(n1291), .C(n24), .D(n1290), .Z(n1006) );
  COND2X1 U997 ( .A(n27), .B(n1292), .C(n24), .D(n1291), .Z(n1007) );
  COND2X1 U998 ( .A(n27), .B(n1293), .C(n24), .D(n1292), .Z(n1008) );
  COND2X1 U999 ( .A(n27), .B(n1294), .C(n24), .D(n1293), .Z(n1009) );
  COND2X1 U1000 ( .A(n27), .B(n1295), .C(n24), .D(n1294), .Z(n1010) );
  COND2X1 U1001 ( .A(n27), .B(n1296), .C(n24), .D(n1295), .Z(n1011) );
  COND2X1 U1002 ( .A(n27), .B(n1297), .C(n24), .D(n1296), .Z(n1012) );
  COND2X1 U1003 ( .A(n27), .B(n1298), .C(n24), .D(n1297), .Z(n1013) );
  COND2X1 U1004 ( .A(n27), .B(n1299), .C(n24), .D(n1298), .Z(n1014) );
  COND2X1 U1005 ( .A(n27), .B(n1300), .C(n24), .D(n1299), .Z(n1015) );
  COND2X1 U1006 ( .A(n27), .B(n1301), .C(n24), .D(n1300), .Z(n1016) );
  COND2X1 U1007 ( .A(n27), .B(n1302), .C(n24), .D(n1301), .Z(n1017) );
  COND2X1 U1008 ( .A(n27), .B(n1303), .C(n24), .D(n1302), .Z(n1018) );
  COND2X1 U1009 ( .A(n27), .B(n1304), .C(n24), .D(n1303), .Z(n1019) );
  COND2X1 U1010 ( .A(n27), .B(n1305), .C(n24), .D(n1304), .Z(n1020) );
  COND2X1 U1011 ( .A(n27), .B(n1306), .C(n24), .D(n1305), .Z(n1021) );
  COND2X1 U1012 ( .A(n27), .B(n1307), .C(n24), .D(n1306), .Z(n1022) );
  COND2X1 U1013 ( .A(n27), .B(n1308), .C(n24), .D(n1307), .Z(n1023) );
  COND2X1 U1014 ( .A(n27), .B(n1309), .C(n24), .D(n1308), .Z(n1024) );
  COND2X1 U1015 ( .A(n27), .B(n1310), .C(n24), .D(n1309), .Z(n1025) );
  COND2X1 U1016 ( .A(n27), .B(n1311), .C(n24), .D(n1310), .Z(n1026) );
  CND2IX1 U1047 ( .B(n1899), .A(n1856), .Z(n1313) );
  COND2X1 U1048 ( .A(n18), .B(n1854), .C(n1344), .D(n15), .Z(n817) );
  COND2X1 U1049 ( .A(n18), .B(n1315), .C(n15), .D(n1314), .Z(n1029) );
  COND2X1 U1052 ( .A(n18), .B(n1318), .C(n15), .D(n1317), .Z(n1032) );
  COND2X1 U1053 ( .A(n18), .B(n1319), .C(n15), .D(n1318), .Z(n1033) );
  COND2X1 U1054 ( .A(n18), .B(n1320), .C(n15), .D(n1319), .Z(n1034) );
  COND2X1 U1055 ( .A(n18), .B(n1321), .C(n15), .D(n1320), .Z(n1035) );
  COND2X1 U1056 ( .A(n18), .B(n1322), .C(n15), .D(n1321), .Z(n1036) );
  COND2X1 U1057 ( .A(n18), .B(n1323), .C(n15), .D(n1322), .Z(n1037) );
  COND2X1 U1058 ( .A(n18), .B(n1324), .C(n15), .D(n1323), .Z(n1038) );
  COND2X1 U1059 ( .A(n18), .B(n1325), .C(n15), .D(n1324), .Z(n1039) );
  COND2X1 U1060 ( .A(n18), .B(n1326), .C(n15), .D(n1325), .Z(n1040) );
  COND2X1 U1061 ( .A(n18), .B(n1327), .C(n15), .D(n1326), .Z(n1041) );
  COND2X1 U1062 ( .A(n18), .B(n1328), .C(n15), .D(n1327), .Z(n1042) );
  COND2X1 U1063 ( .A(n18), .B(n1329), .C(n15), .D(n1328), .Z(n1043) );
  COND2X1 U1064 ( .A(n18), .B(n1330), .C(n15), .D(n1329), .Z(n1044) );
  COND2X1 U1065 ( .A(n18), .B(n1331), .C(n15), .D(n1330), .Z(n1045) );
  COND2X1 U1066 ( .A(n18), .B(n1332), .C(n15), .D(n1331), .Z(n1046) );
  COND2X1 U1067 ( .A(n18), .B(n1333), .C(n15), .D(n1332), .Z(n1047) );
  COND2X1 U1068 ( .A(n18), .B(n1334), .C(n15), .D(n1333), .Z(n1048) );
  COND2X1 U1069 ( .A(n18), .B(n1335), .C(n15), .D(n1334), .Z(n1049) );
  COND2X1 U1070 ( .A(n18), .B(n1336), .C(n15), .D(n1335), .Z(n1050) );
  COND2X1 U1071 ( .A(n18), .B(n1337), .C(n15), .D(n1336), .Z(n1051) );
  COND2X1 U1072 ( .A(n18), .B(n1338), .C(n15), .D(n1337), .Z(n1052) );
  COND2X1 U1073 ( .A(n18), .B(n1339), .C(n15), .D(n1338), .Z(n1053) );
  COND2X1 U1075 ( .A(n18), .B(n1341), .C(n15), .D(n1340), .Z(n1055) );
  CND2IX1 U1109 ( .B(n1899), .A(n1850), .Z(n1344) );
  CENX2 U1244 ( .A(n1878), .B(a[16]), .Z(n74) );
  CENX2 U1253 ( .A(n1869), .B(a[10]), .Z(n50) );
  CFD1QXL clk_r_REG173_S1 ( .D(n376), .CP(n1823), .Q(n1815) );
  CFD1QXL clk_r_REG116_S1 ( .D(n378), .CP(n1823), .Q(n1813) );
  CFD1QXL clk_r_REG170_S1 ( .D(n380), .CP(n1823), .Q(n1811) );
  CFD1QXL clk_r_REG171_S1 ( .D(n381), .CP(n1823), .Q(n1810) );
  CFD1QXL clk_r_REG26_S1 ( .D(n379), .CP(n1823), .Q(n1812) );
  CFD1QXL clk_r_REG2_S1 ( .D(n399), .CP(n1823), .Q(n1792) );
  CFD1QXL clk_r_REG127_S1 ( .D(n401), .CP(n1823), .Q(n1790) );
  CFD1QXL clk_r_REG42_S1 ( .D(n760), .CP(n1823), .Q(n1657) );
  CFD1QXL clk_r_REG107_S1 ( .D(n458), .CP(n1823), .Q(n1770) );
  CFD1QXL clk_r_REG99_S1 ( .D(n578), .CP(n1823), .Q(n1723) );
  CFD1QXL clk_r_REG62_S1 ( .D(n573), .CP(n1823), .Q(n1728) );
  CFD1QXL clk_r_REG174_S1 ( .D(n436), .CP(n1823), .Q(n1774) );
  CFD1QXL clk_r_REG56_S1 ( .D(n459), .CP(n1823), .Q(n1769) );
  CFD1QXL clk_r_REG137_S1 ( .D(n783), .CP(n1823), .Q(n1648) );
  CFD1QXL clk_r_REG74_S1 ( .D(n530), .CP(n1823), .Q(n1743) );
  CFD1QXL clk_r_REG72_S1 ( .D(n506), .CP(n1823), .Q(n1752) );
  CFD1QXL clk_r_REG38_S1 ( .D(n616), .CP(n1823), .Q(n1711) );
  CFD1QXL clk_r_REG12_S1 ( .D(n714), .CP(n1823), .Q(n1675) );
  CFD1QXL clk_r_REG25_S1 ( .D(n770), .CP(n1823), .Q(n1653) );
  CFD1QXL clk_r_REG189_S1 ( .D(n536), .CP(n1823), .Q(n1737) );
  CFD1QXL clk_r_REG78_S1 ( .D(n620), .CP(n1823), .Q(n1707) );
  CFD1QXL clk_r_REG142_S1 ( .D(n794), .CP(n1823), .Q(n1643) );
  CFD1QXL clk_r_REG36_S1 ( .D(n600), .CP(n1823), .Q(n1715) );
  CFD1QXL clk_r_REG14_S1 ( .D(n700), .CP(n1823), .Q(n1681) );
  CFD1QXL clk_r_REG41_S1 ( .D(n759), .CP(n1823), .Q(n1658) );
  CFD1QXL clk_r_REG157_S1 ( .D(n749), .CP(n1823), .Q(n1662) );
  CFD1QXL clk_r_REG8_S1 ( .D(n480), .CP(n1823), .Q(n1762) );
  CFD1QXL clk_r_REG4_S1 ( .D(n377), .CP(n1823), .Q(n1814) );
  CFD1QXL clk_r_REG27_S1 ( .D(n403), .CP(n1823), .Q(n1788) );
  CFD1QXL clk_r_REG114_S1 ( .D(n405), .CP(n1823), .Q(n1786) );
  CFD1QXL clk_r_REG146_S1 ( .D(n319), .CP(n1823), .Q(n1821) );
  CFD1QXL clk_r_REG150_S1 ( .D(n327), .CP(n1823), .Q(n1818) );
  CFD1QXL clk_r_REG148_S1 ( .D(n1624), .CP(n1823), .Q(n1822) );
  CFD1QXL clk_r_REG145_S1 ( .D(n320), .CP(n1823), .Q(n1820) );
  CFD1QXL clk_r_REG149_S1 ( .D(n328), .CP(n1823), .Q(n1817) );
  CFD1QXL clk_r_REG7_S1 ( .D(n479), .CP(n1823), .Q(n1763) );
  CFD1QXL clk_r_REG135_S1 ( .D(n767), .CP(n1823), .Q(n1656) );
  CFD1QXL clk_r_REG124_S1 ( .D(n726), .CP(n1823), .Q(n1671) );
  CFD1QXL clk_r_REG82_S1 ( .D(n580), .CP(n1823), .Q(n1721) );
  CFD1QXL clk_r_REG63_S1 ( .D(n574), .CP(n1823), .Q(n1727) );
  CFD1QXL clk_r_REG34_S1 ( .D(n556), .CP(n1823), .Q(n1733) );
  CFD1QXL clk_r_REG95_S1 ( .D(n686), .CP(n1823), .Q(n1685) );
  CFD1QXL clk_r_REG1_S1 ( .D(n778), .CP(n1823), .Q(n1795) );
  CFD1QXL clk_r_REG105_S1 ( .D(n532), .CP(n1823), .Q(n1741) );
  CFD1QXL clk_r_REG111_S1 ( .D(n508), .CP(n1823), .Q(n1750) );
  CFD1QXL clk_r_REG88_S1 ( .D(n618), .CP(n1823), .Q(n1709) );
  CFD1QXL clk_r_REG158_S1 ( .D(n750), .CP(n1823), .Q(n1661) );
  CFD1QXL clk_r_REG3_S1 ( .D(n400), .CP(n1823), .Q(n1791) );
  CFD1QXL clk_r_REG28_S1 ( .D(n404), .CP(n1823), .Q(n1787) );
  CFD1QXL clk_r_REG130_S1 ( .D(n482), .CP(n1823), .Q(n1760) );
  CFD1QXL clk_r_REG138_S1 ( .D(n784), .CP(n1823), .Q(n1647) );
  CFD1QXL clk_r_REG143_S1 ( .D(n797), .CP(n1823), .Q(n1793) );
  CFD1QXL clk_r_REG69_S1 ( .D(n596), .CP(n1823), .Q(n1719) );
  CFD1QXL clk_r_REG141_S1 ( .D(n793), .CP(n1823), .Q(n1644) );
  CFD1QXL clk_r_REG18_S1 ( .D(n738), .CP(n1823), .Q(n1665) );
  CFD1QXL clk_r_REG123_S1 ( .D(n725), .CP(n1823), .Q(n1672) );
  CFD1QXL clk_r_REG122_S1 ( .D(n740), .CP(n1823), .Q(n1663) );
  CFD1QXL clk_r_REG40_S1 ( .D(n634), .CP(n1823), .Q(n1705) );
  CFD1QXL clk_r_REG24_S1 ( .D(n769), .CP(n1823), .Q(n1654) );
  CFD1QXL clk_r_REG187_S1 ( .D(n462), .CP(n1823), .Q(n1766) );
  CFD1QXL clk_r_REG100_S1 ( .D(n597), .CP(n1823), .Q(n1718) );
  CFD1QXL clk_r_REG165_S1 ( .D(n434), .CP(n1823), .Q(n1775) );
  CFD1QXL clk_r_REG16_S1 ( .D(n728), .CP(n1823), .Q(n1669) );
  CFD1QXL clk_r_REG103_S1 ( .D(n558), .CP(n1823), .Q(n1731) );
  CFD1QXL clk_r_REG49_S1 ( .D(n688), .CP(n1823), .Q(n1683) );
  CFD1QXL clk_r_REG32_S1 ( .D(n534), .CP(n1823), .Q(n1739) );
  CFD1QXL clk_r_REG169_S1 ( .D(n997), .CP(n1823), .Q(n1635) );
  CFD1QXL clk_r_REG59_S1 ( .D(n484), .CP(n1823), .Q(n1758) );
  CFD1QXL clk_r_REG139_S1 ( .D(n787), .CP(n1823), .Q(n1646) );
  CFD1QXL clk_r_REG53_S1 ( .D(n652), .CP(n1823), .Q(n1697) );
  CFD1QXL clk_r_REG20_S1 ( .D(n752), .CP(n1823), .Q(n1659) );
  CFD1QXL clk_r_REG156_S1 ( .D(n790), .CP(n1823), .Q(n1794) );
  CFD1QXL clk_r_REG167_S1 ( .D(n1026), .CP(n1823), .Q(n1634) );
  CFD1QXL clk_r_REG51_S1 ( .D(n670), .CP(n1823), .Q(n1691) );
  CFD1QXL clk_r_REG154_S1 ( .D(n781), .CP(n1823), .Q(n1650) );
  CFD1QXL clk_r_REG118_S1 ( .D(n329), .CP(n1823), .Q(n1816) );
  CFD1QX2 clk_r_REG70_S1 ( .D(n958), .CP(n1823), .Q(n1639) );
  CFD1QX1 clk_r_REG185_S1 ( .D(n581), .CP(n1823), .Q(n1807) );
  CFD1QX2 clk_r_REG81_S1 ( .D(n579), .CP(n1823), .Q(n1722) );
  CFD1QX2 clk_r_REG109_S1 ( .D(n430), .CP(n1823), .Q(n1779) );
  CFD1QX2 clk_r_REG134_S1 ( .D(n576), .CP(n1823), .Q(n1725) );
  CFD1QX2 clk_r_REG30_S1 ( .D(n432), .CP(n1823), .Q(n1777) );
  CFD1QX2 clk_r_REG190_S1 ( .D(n601), .CP(n1823), .Q(n1714) );
  CFD1QX1 clk_r_REG166_S1 ( .D(n923), .CP(n1823), .Q(n1641) );
  CFD1QX1 clk_r_REG188_S1 ( .D(n535), .CP(n1823), .Q(n1738) );
  CFD1QX1 clk_r_REG35_S1 ( .D(n599), .CP(n1823), .Q(n1716) );
  CFD1QX2 clk_r_REG168_S1 ( .D(n995), .CP(n1823), .Q(n1631) );
  CFD1QX2 clk_r_REG128_S1 ( .D(n402), .CP(n1823), .Q(n1789) );
  CFD1QX1 clk_r_REG151_S1 ( .D(n1073), .CP(n1823), .Q(n1633) );
  CFD1QX2 clk_r_REG181_S1 ( .D(n538), .CP(n1823), .Q(n1808) );
  CFD1QX2 clk_r_REG11_S1 ( .D(n713), .CP(n1823), .Q(n1676) );
  CFD1QX2 clk_r_REG96_S1 ( .D(n715), .CP(n1823), .Q(n1674) );
  CFD1QX1 clk_r_REG66_S1 ( .D(n964), .CP(n1823), .Q(n1637) );
  CFD1QX1 clk_r_REG64_S1 ( .D(n689), .CP(n1823), .Q(n1803) );
  CFD1QX1 clk_r_REG31_S1 ( .D(n533), .CP(n1823), .Q(n1740) );
  CFD1QX1 clk_r_REG91_S1 ( .D(n658), .CP(n1823), .Q(n1804) );
  CFD1QX1 clk_r_REG83_S1 ( .D(n673), .CP(n1823), .Q(n1688) );
  CFD1QX1 clk_r_REG112_S1 ( .D(n485), .CP(n1823), .Q(n1757) );
  CFD1QX1 clk_r_REG75_S1 ( .D(n703), .CP(n1823), .Q(n1678) );
  CFD1QX1 clk_r_REG46_S1 ( .D(n701), .CP(n1823), .Q(n1680) );
  CFD1QX2 clk_r_REG58_S1 ( .D(n483), .CP(n1823), .Q(n1759) );
  CFD1QX1 clk_r_REG176_S1 ( .D(n464), .CP(n1823), .Q(n1764) );
  CFD1QX1 clk_r_REG86_S1 ( .D(n640), .CP(n1823), .Q(n1699) );
  CFD1QX1 clk_r_REG60_S1 ( .D(n509), .CP(n1823), .Q(n1749) );
  CFD1QX2 clk_r_REG73_S1 ( .D(n529), .CP(n1823), .Q(n1744) );
  CFD1QX1 clk_r_REG37_S1 ( .D(n615), .CP(n1823), .Q(n1712) );
  CFD1QX1 clk_r_REG192_S1 ( .D(n621), .CP(n1823), .Q(n1806) );
  CFD1QX1 clk_r_REG65_S1 ( .D(n690), .CP(n1823), .Q(n1802) );
  CFD1QX2 clk_r_REG104_S1 ( .D(n531), .CP(n1823), .Q(n1742) );
  CFD1QX1 clk_r_REG45_S1 ( .D(n945), .CP(n1823), .Q(n1640) );
  CFD1QX2 clk_r_REG101_S1 ( .D(n598), .CP(n1823), .Q(n1717) );
  CFD1QX1 clk_r_REG110_S1 ( .D(n507), .CP(n1823), .Q(n1751) );
  CFD1QX1 clk_r_REG183_S1 ( .D(n559), .CP(n1823), .Q(n1730) );
  CFD1QX1 clk_r_REG159_S1 ( .D(n742), .CP(n1823), .Q(n1799) );
  CFD1QX1 clk_r_REG191_S1 ( .D(n602), .CP(n1823), .Q(n1713) );
  CFD1QX1 clk_r_REG90_S1 ( .D(n638), .CP(n1823), .Q(n1701) );
  CFD1QX1 clk_r_REG153_S1 ( .D(n636), .CP(n1823), .Q(n1703) );
  CFD1QX1 clk_r_REG77_S1 ( .D(n619), .CP(n1823), .Q(n1708) );
  CFD1QX1 clk_r_REG180_S1 ( .D(n514), .CP(n1823), .Q(n1745) );
  CFD1QX1 clk_r_REG93_S1 ( .D(n718), .CP(n1823), .Q(n1800) );
  CFD1QX1 clk_r_REG125_S1 ( .D(n653), .CP(n1823), .Q(n1696) );
  CFD1QX1 clk_r_REG129_S1 ( .D(n481), .CP(n1823), .Q(n1761) );
  CFD1QX1 clk_r_REG164_S1 ( .D(n433), .CP(n1823), .Q(n1776) );
  CFD1QX2 clk_r_REG98_S1 ( .D(n577), .CP(n1823), .Q(n1724) );
  CFD1QX2 clk_r_REG68_S1 ( .D(n595), .CP(n1823), .Q(n1720) );
  CFD1QX2 clk_r_REG113_S1 ( .D(n486), .CP(n1823), .Q(n1756) );
  CFD1QX2 clk_r_REG71_S1 ( .D(n505), .CP(n1823), .Q(n1753) );
  CFD1QX2 clk_r_REG179_S1 ( .D(n488), .CP(n1823), .Q(n1754) );
  CFD1QX2 clk_r_REG160_S1 ( .D(n671), .CP(n1823), .Q(n1690) );
  CFD1QX1 clk_r_REG175_S1 ( .D(n463), .CP(n1823), .Q(n1765) );
  CFD1QX1 clk_r_REG0_S1 ( .D(n777), .CP(n1823), .Q(n1796) );
  CFD1QX1 clk_r_REG22_S1 ( .D(n775), .CP(n1823), .Q(n1652) );
  CFD1QX1 clk_r_REG55_S1 ( .D(n762), .CP(n1823), .Q(n1797) );
  CFD1QX1 clk_r_REG29_S1 ( .D(n431), .CP(n1823), .Q(n1778) );
  CFD1QX1 clk_r_REG102_S1 ( .D(n557), .CP(n1823), .Q(n1732) );
  CFD1QX1 clk_r_REG172_S1 ( .D(n410), .CP(n1823), .Q(n1783) );
  CFD1QX1 clk_r_REG133_S1 ( .D(n575), .CP(n1823), .Q(n1726) );
  CFD1QX2 clk_r_REG80_S1 ( .D(n656), .CP(n1823), .Q(n1693) );
  CFD1QX2 clk_r_REG126_S1 ( .D(n654), .CP(n1823), .Q(n1695) );
  CFD1QX1 clk_r_REG13_S1 ( .D(n699), .CP(n1823), .Q(n1682) );
  CFD1QX2 clk_r_REG43_S1 ( .D(n729), .CP(n1823), .Q(n1668) );
  CFD1QX2 clk_r_REG94_S1 ( .D(n685), .CP(n1823), .Q(n1686) );
  CFD1QX1 clk_r_REG17_S1 ( .D(n737), .CP(n1823), .Q(n1666) );
  CFD1QX1 clk_r_REG9_S1 ( .D(n455), .CP(n1823), .Q(n1773) );
  CFD1QX1 clk_r_REG50_S1 ( .D(n669), .CP(n1823), .Q(n1692) );
  CFD1QX1 clk_r_REG186_S1 ( .D(n461), .CP(n1823), .Q(n1767) );
  CFD1QX2 clk_r_REG163_S1 ( .D(n512), .CP(n1823), .Q(n1746) );
  CFD1QX1 clk_r_REG182_S1 ( .D(n408), .CP(n1823), .Q(n1784) );
  CFD1QX1 clk_r_REG84_S1 ( .D(n674), .CP(n1823), .Q(n1687) );
  CFD1QX1 clk_r_REG121_S1 ( .D(n739), .CP(n1823), .Q(n1664) );
  CFD1QX1 clk_r_REG44_S1 ( .D(n730), .CP(n1823), .Q(n1667) );
  CFD1QX1 clk_r_REG87_S1 ( .D(n617), .CP(n1823), .Q(n1710) );
  CFD1QX1 clk_r_REG33_S1 ( .D(n555), .CP(n1823), .Q(n1734) );
  CFD1QX1 clk_r_REG120_S1 ( .D(n1078), .CP(n1823), .Q(n1632) );
  CFD1QXL clk_r_REG140_S1 ( .D(n788), .CP(n1823), .Q(n1645) );
  CFD1QXL clk_r_REG23_S1 ( .D(n776), .CP(n1823), .Q(n1651) );
  CFD1QXL clk_r_REG155_S1 ( .D(n782), .CP(n1823), .Q(n1649) );
  CFD1QXL clk_r_REG136_S1 ( .D(n768), .CP(n1823), .Q(n1655) );
  CFD1QXL clk_r_REG147_S1 ( .D(n325), .CP(n1823), .Q(n1819) );
  CFD1QXL clk_r_REG144_S1 ( .D(n795), .CP(n1823), .Q(n1642) );
  CFD1QX1 clk_r_REG108_S1 ( .D(n429), .CP(n1823), .Q(n1780) );
  CFD1QX1 clk_r_REG10_S1 ( .D(n456), .CP(n1823), .Q(n1772) );
  CFD1QX2 clk_r_REG89_S1 ( .D(n637), .CP(n1823), .Q(n1702) );
  CFD1QX1 clk_r_REG131_S1 ( .D(n553), .CP(n1823), .Q(n1736) );
  CFD1QX1 clk_r_REG54_S1 ( .D(n761), .CP(n1823), .Q(n1798) );
  CFD1QX2 clk_r_REG61_S1 ( .D(n510), .CP(n1823), .Q(n1748) );
  CFD1QX2 clk_r_REG57_S1 ( .D(n460), .CP(n1823), .Q(n1768) );
  CFD1QX2 clk_r_REG67_S1 ( .D(n961), .CP(n1823), .Q(n1638) );
  CFD1QX2 clk_r_REG21_S1 ( .D(n971), .CP(n1823), .Q(n1636) );
  CFD1QX1 clk_r_REG6_S1 ( .D(n428), .CP(n1823), .Q(n1781) );
  CFD1QX1 clk_r_REG48_S1 ( .D(n687), .CP(n1823), .Q(n1684) );
  CFD1QX4 clk_r_REG92_S1 ( .D(n717), .CP(n1823), .Q(n1801) );
  CFD1QX1 clk_r_REG76_S1 ( .D(n704), .CP(n1823), .Q(n1677) );
  CFD1QX1 clk_r_REG106_S1 ( .D(n457), .CP(n1823), .Q(n1771) );
  CFD1QX2 clk_r_REG178_S1 ( .D(n487), .CP(n1823), .Q(n1755) );
  CFD1QX4 clk_r_REG177_S1 ( .D(n489), .CP(n1823), .Q(n1809) );
  CFD1QX1 clk_r_REG152_S1 ( .D(n635), .CP(n1823), .Q(n1704) );
  CFD1QX1 clk_r_REG47_S1 ( .D(n702), .CP(n1823), .Q(n1679) );
  CFD1QX1 clk_r_REG5_S1 ( .D(n427), .CP(n1823), .Q(n1782) );
  CFD1QX2 clk_r_REG19_S1 ( .D(n751), .CP(n1823), .Q(n1660) );
  CFD1QX1 clk_r_REG184_S1 ( .D(n560), .CP(n1823), .Q(n1729) );
  CFD1QX2 clk_r_REG161_S1 ( .D(n672), .CP(n1823), .Q(n1689) );
  CFD1QX2 clk_r_REG15_S1 ( .D(n727), .CP(n1823), .Q(n1670) );
  CFD1QX4 clk_r_REG162_S1 ( .D(n511), .CP(n1823), .Q(n1747) );
  CFD1QX2 clk_r_REG132_S1 ( .D(n554), .CP(n1823), .Q(n1735) );
  CFD1QX1 clk_r_REG97_S1 ( .D(n716), .CP(n1823), .Q(n1673) );
  CFD1QX2 clk_r_REG79_S1 ( .D(n655), .CP(n1823), .Q(n1694) );
  CFD1QX1 clk_r_REG39_S1 ( .D(n633), .CP(n1823), .Q(n1706) );
  CFD1QX4 clk_r_REG85_S1 ( .D(n639), .CP(n1823), .Q(n1700) );
  CFD1QX4 clk_r_REG193_S1 ( .D(n622), .CP(n1823), .Q(n1805) );
  CFD1QX2 clk_r_REG115_S1 ( .D(n406), .CP(n1823), .Q(n1785) );
  CFD1QX2 clk_r_REG52_S1 ( .D(n651), .CP(n1823), .Q(n1698) );
  COND2X1 U1131 ( .A(1'b1), .B(n1366), .C(n6), .D(n1365), .Z(n1079) );
  COND2X1 U1118 ( .A(1'b1), .B(n1353), .C(n6), .D(n1352), .Z(n1066) );
  COND2X1 U1117 ( .A(1'b1), .B(n1352), .C(n6), .D(n1351), .Z(n1065) );
  COND2X1 U1114 ( .A(1'b1), .B(n1349), .C(n6), .D(n1348), .Z(n1062) );
  CNR2X2 U1271 ( .A(n6), .B(n1366), .Z(n1080) );
  CNR2X2 U1272 ( .A(n6), .B(n1367), .Z(n1081) );
  CNR2X2 U1273 ( .A(n6), .B(n1368), .Z(n1082) );
  CNR2X2 U1274 ( .A(n6), .B(n1369), .Z(n1083) );
  CNR2X2 U1275 ( .A(n6), .B(n1370), .Z(n1084) );
  CNR2X2 U1276 ( .A(n6), .B(n1371), .Z(n1085) );
  CNR2X2 U1277 ( .A(n6), .B(n1372), .Z(n1086) );
  CNR2X2 U1278 ( .A(n6), .B(n1373), .Z(n1087) );
  CNR2X2 U1279 ( .A(n6), .B(n1375), .Z(n1089) );
  CNR2X2 U1280 ( .A(n6), .B(n1363), .Z(n1077) );
  CNR2X2 U1281 ( .A(n6), .B(n1362), .Z(n1076) );
  CNR2X2 U1282 ( .A(n6), .B(n1361), .Z(n1075) );
  CNR2X2 U1283 ( .A(n6), .B(n1360), .Z(n1074) );
  CNR2X2 U1284 ( .A(n6), .B(n1359), .Z(n1073) );
  CNR2X2 U1285 ( .A(n6), .B(n1358), .Z(n1072) );
  CNR2X2 U1286 ( .A(n6), .B(n1357), .Z(n1071) );
  CNR2X2 U1287 ( .A(n6), .B(n1356), .Z(n1070) );
  CNR2X2 U1288 ( .A(n6), .B(n1355), .Z(n1069) );
  CNR2X2 U1289 ( .A(n6), .B(n1354), .Z(n1068) );
  CNR2X2 U1290 ( .A(n6), .B(n1364), .Z(n1078) );
  CNR2X2 U1291 ( .A(n6), .B(n1374), .Z(n1088) );
  CNR2X2 U1292 ( .A(n6), .B(n1350), .Z(n1064) );
  CNR2X2 U1293 ( .A(n6), .B(n1353), .Z(n1067) );
  CNR2X2 U1294 ( .A(n6), .B(n1349), .Z(n1063) );
  CNR2X2 U1295 ( .A(n6), .B(n1345), .Z(n1059) );
  CNR2X2 U1296 ( .A(n6), .B(n1347), .Z(n1061) );
  CNR2X2 U1297 ( .A(n6), .B(n1346), .Z(n1060) );
  CIVX2 U1298 ( .A(n1393), .Z(n1360) );
  CIVX2 U1299 ( .A(n1846), .Z(n1364) );
  CIVX2 U1300 ( .A(n1849), .Z(n1361) );
  CIVX2 U1301 ( .A(n1847), .Z(n1363) );
  CIVX2 U1302 ( .A(n1550), .Z(n1358) );
  CIVX2 U1303 ( .A(n1848), .Z(n1362) );
  CIVX2 U1304 ( .A(n1392), .Z(n1359) );
  CIVX2 U1305 ( .A(n1089), .Z(n335) );
  CIVX2 U1306 ( .A(n335), .Z(product[1]) );
  CIVX2 U1307 ( .A(n1842), .Z(n1368) );
  CIVX2 U1308 ( .A(n1840), .Z(n1370) );
  CIVX2 U1309 ( .A(n1845), .Z(n1365) );
  CIVX2 U1310 ( .A(n1839), .Z(n1371) );
  CIVX2 U1311 ( .A(n1844), .Z(n1366) );
  CIVX2 U1312 ( .A(n1843), .Z(n1367) );
  CIVX2 U1313 ( .A(n1837), .Z(n1373) );
  CIVX2 U1314 ( .A(n1838), .Z(n1372) );
  CIVX2 U1315 ( .A(n1407), .Z(n1374) );
  CIVX2 U1316 ( .A(n1408), .Z(n1375) );
  CIVX2 U1317 ( .A(a[2]), .Z(n15) );
  CIVX2 U1318 ( .A(b[31]), .Z(n1345) );
  CIVX2 U1319 ( .A(n331), .Z(n329) );
  CIVX2 U1320 ( .A(n148), .Z(product[2]) );
  CIVX2 U1321 ( .A(n1554), .Z(n1357) );
  CIVX2 U1322 ( .A(n1841), .Z(n1369) );
  CIVX2 U1323 ( .A(b[25]), .Z(n1351) );
  CIVX2 U1324 ( .A(b[24]), .Z(n1352) );
  CIVX2 U1325 ( .A(n1389), .Z(n1356) );
  CIVX2 U1326 ( .A(n1387), .Z(n1354) );
  CIVX2 U1327 ( .A(b[26]), .Z(n1350) );
  CIVX2 U1328 ( .A(n1386), .Z(n1353) );
  CIVX2 U1329 ( .A(b[30]), .Z(n1346) );
  CIVX2 U1330 ( .A(b[28]), .Z(n1348) );
  CIVX2 U1331 ( .A(b[27]), .Z(n1349) );
  CIVX2 U1332 ( .A(b[29]), .Z(n1347) );
  CIVX2 U1333 ( .A(n1388), .Z(n1355) );
  CIVXL U1335 ( .A(n195), .Z(n1548) );
  CIVX2 U1336 ( .A(n1391), .Z(n1549) );
  CIVX4 U1337 ( .A(n1549), .Z(n1550) );
  CANR1X1 U1338 ( .A(n343), .B(n194), .C(n191), .Z(n189) );
  CANR1XL U1339 ( .A(n181), .B(n194), .C(n1561), .Z(n180) );
  CENXL U1340 ( .A(n1862), .B(n1388), .Z(n1262) );
  CENXL U1341 ( .A(n1867), .B(n1388), .Z(n1235) );
  CENXL U1342 ( .A(n1851), .B(n1388), .Z(n1322) );
  CENXL U1343 ( .A(n1855), .B(n1388), .Z(n1291) );
  CENXL U1344 ( .A(n1872), .B(n1388), .Z(n1210) );
  COR2X1 U1345 ( .A(n584), .B(n603), .Z(n1551) );
  CENX1 U1346 ( .A(n1562), .B(n1638), .Z(n614) );
  CEO3XL U1347 ( .A(n909), .B(n951), .C(n1059), .Z(n377) );
  CND2XL U1348 ( .A(n1551), .B(n223), .Z(n128) );
  CIVX2 U1349 ( .A(n546), .Z(n1581) );
  CIVX2 U1350 ( .A(n1390), .Z(n1552) );
  CIVXL U1351 ( .A(n1552), .Z(n1553) );
  CIVX1 U1352 ( .A(n1552), .Z(n1554) );
  CIVX2 U1353 ( .A(n1552), .Z(n1555) );
  CANR1X1 U1354 ( .A(n228), .B(n1612), .C(n221), .Z(n1556) );
  CANR1X1 U1355 ( .A(n228), .B(n1612), .C(n221), .Z(n215) );
  CFA1XL U1356 ( .A(n968), .B(n1018), .CI(n1046), .CO(n727), .S(n728) );
  CFA1X1 U1357 ( .A(n922), .B(n1042), .CI(n1014), .CO(n671), .S(n672) );
  COND1X2 U1358 ( .A(n193), .B(n187), .C(n188), .Z(n182) );
  CNR2X1 U1359 ( .A(n248), .B(n251), .Z(n246) );
  CNR2X2 U1360 ( .A(n660), .B(n675), .Z(n248) );
  CFA1XL U1361 ( .A(n928), .B(n970), .CI(n948), .CO(n751), .S(n752) );
  COND1X1 U1362 ( .A(n167), .B(n195), .C(n168), .Z(n166) );
  CAN2X1 U1363 ( .A(n1613), .B(n1614), .Z(n1609) );
  CANR1X2 U1364 ( .A(n261), .B(n1617), .C(n254), .Z(n252) );
  CENX1 U1365 ( .A(n1850), .B(b[27]), .Z(n1316) );
  CND2XL U1366 ( .A(n1735), .B(n571), .Z(n1591) );
  CND2XL U1367 ( .A(n552), .B(n571), .Z(n1592) );
  CENX1 U1368 ( .A(n1886), .B(a[20]), .Z(n89) );
  CIVX2 U1369 ( .A(n1865), .Z(n1861) );
  CIVX1 U1370 ( .A(n1854), .Z(n1851) );
  CIVX2 U1371 ( .A(n39), .Z(n1871) );
  CIVX1 U1372 ( .A(n12), .Z(n1854) );
  COND2X2 U1373 ( .A(n36), .B(n1266), .C(n1265), .D(n1606), .Z(n982) );
  COND2X2 U1374 ( .A(n36), .B(n1260), .C(n1259), .D(n1606), .Z(n976) );
  COND2X2 U1375 ( .A(n53), .B(n1212), .C(n1211), .D(n50), .Z(n930) );
  CEOXL U1376 ( .A(a[6]), .B(n1861), .Z(n1422) );
  CENX2 U1377 ( .A(n1857), .B(a[6]), .Z(n1606) );
  CIVXL U1378 ( .A(n113), .Z(n1435) );
  COND2X1 U1379 ( .A(n53), .B(n1216), .C(n1215), .D(n50), .Z(n934) );
  CIVXL U1380 ( .A(n265), .Z(n264) );
  COND2X2 U1381 ( .A(n27), .B(n1602), .C(n1285), .D(n24), .Z(n1001) );
  CENX1 U1382 ( .A(n1858), .B(b[27]), .Z(n1285) );
  CENXL U1383 ( .A(n1557), .B(n180), .Z(product[27]) );
  CAN2XL U1384 ( .A(n341), .B(n179), .Z(n1557) );
  CANR1X1 U1385 ( .A(n210), .B(n1621), .C(n201), .Z(n199) );
  CENXL U1386 ( .A(n1558), .B(n152), .Z(product[31]) );
  CAN2X1 U1387 ( .A(n1623), .B(n151), .Z(n1558) );
  CNIVX1 U1388 ( .A(n1901), .Z(product[3]) );
  CNIVX1 U1389 ( .A(n1900), .Z(product[5]) );
  COND1X2 U1390 ( .A(n281), .B(n275), .C(n276), .Z(n274) );
  CEO3XL U1391 ( .A(n875), .B(n929), .C(n1001), .Z(n379) );
  COND2X2 U1392 ( .A(n18), .B(n1317), .C(n1316), .D(n15), .Z(n1031) );
  CANR1X1 U1393 ( .A(n169), .B(n182), .C(n170), .Z(n168) );
  CIVX1 U1394 ( .A(n182), .Z(n184) );
  COND1X1 U1395 ( .A(n1600), .B(n215), .C(n199), .Z(n197) );
  CENXL U1396 ( .A(n1850), .B(b[28]), .Z(n1315) );
  CANR1X2 U1397 ( .A(n241), .B(n1618), .C(n236), .Z(n234) );
  CIVXL U1398 ( .A(n184), .Z(n1561) );
  CENX2 U1399 ( .A(n1700), .B(n1805), .Z(n1562) );
  CFA1XL U1400 ( .A(n854), .B(n914), .CI(n866), .CO(n511), .S(n512) );
  CIVXL U1401 ( .A(n187), .Z(n342) );
  CFA1XL U1402 ( .A(n905), .B(n1015), .CI(n989), .CO(n685), .S(n686) );
  CFA1XL U1403 ( .A(n908), .B(n946), .CI(n926), .CO(n729), .S(n730) );
  COND2XL U1404 ( .A(n61), .B(n1204), .C(n1203), .D(n58), .Z(n923) );
  COND2XL U1405 ( .A(n61), .B(n1195), .C(n1194), .D(n58), .Z(n914) );
  COND2XL U1406 ( .A(n61), .B(n1205), .C(n1204), .D(n58), .Z(n924) );
  COND2XL U1407 ( .A(n61), .B(n1200), .C(n1199), .D(n58), .Z(n919) );
  COND2XL U1408 ( .A(n61), .B(n1201), .C(n1200), .D(n58), .Z(n920) );
  COND2XL U1409 ( .A(n61), .B(n1207), .C(n1206), .D(n58), .Z(n926) );
  COND2XL U1410 ( .A(n61), .B(n1203), .C(n1202), .D(n58), .Z(n922) );
  CND2X4 U1411 ( .A(n1605), .B(n58), .Z(n61) );
  CENXL U1412 ( .A(n213), .B(n127), .Z(product[23]) );
  CENXL U1413 ( .A(n1563), .B(n161), .Z(product[30]) );
  CAN2XL U1414 ( .A(n1613), .B(n160), .Z(n1563) );
  CNIVX3 U1415 ( .A(n1395), .Z(n1848) );
  COND2X1 U1416 ( .A(n77), .B(n1155), .C(n1154), .D(n74), .Z(n876) );
  COND1XL U1417 ( .A(n290), .B(n286), .C(n287), .Z(n285) );
  CANR1X2 U1418 ( .A(n1620), .B(n274), .C(n269), .Z(n267) );
  CANR1X1 U1419 ( .A(n301), .B(n1626), .C(n296), .Z(n294) );
  CND2X1 U1420 ( .A(n1626), .B(n1625), .Z(n293) );
  CANR1X1 U1421 ( .A(n1627), .B(n310), .C(n307), .Z(n305) );
  CEO3X1 U1422 ( .A(n1717), .B(n613), .C(n1719), .Z(n590) );
  CND2X1 U1423 ( .A(n1717), .B(n613), .Z(n1564) );
  CND2X1 U1424 ( .A(n1717), .B(n1719), .Z(n1565) );
  CND2X1 U1425 ( .A(n613), .B(n1719), .Z(n1566) );
  CND3X2 U1426 ( .A(n1564), .B(n1565), .C(n1566), .Z(n589) );
  CEOXL U1427 ( .A(n591), .B(n572), .Z(n1567) );
  CEOX1 U1428 ( .A(n1567), .B(n589), .Z(n566) );
  CND2X1 U1429 ( .A(n591), .B(n572), .Z(n1568) );
  CND2X1 U1430 ( .A(n591), .B(n589), .Z(n1569) );
  CND2X1 U1431 ( .A(n572), .B(n589), .Z(n1570) );
  CND3X2 U1432 ( .A(n1568), .B(n1569), .C(n1570), .Z(n565) );
  CND2X1 U1433 ( .A(n1621), .B(n1611), .Z(n1600) );
  CFA1XL U1434 ( .A(n899), .B(n1037), .CI(n983), .CO(n577), .S(n578) );
  CENXL U1435 ( .A(n104), .B(a[28]), .Z(n110) );
  CENXL U1436 ( .A(n104), .B(n1838), .Z(n1099) );
  CENXL U1437 ( .A(n104), .B(n1837), .Z(n1100) );
  CND2XL U1438 ( .A(n104), .B(n1407), .Z(n1825) );
  CND2IXL U1439 ( .B(n1899), .A(n104), .Z(n1104) );
  CENXL U1440 ( .A(n104), .B(n1839), .Z(n1098) );
  CENXL U1441 ( .A(n104), .B(n1408), .Z(n1102) );
  CENXL U1442 ( .A(n1898), .B(n104), .Z(n1103) );
  CND2IX1 U1443 ( .B(n567), .A(n565), .Z(n1585) );
  CENXL U1444 ( .A(n109), .B(n1837), .Z(n1093) );
  CND2IXL U1445 ( .B(n1899), .A(n109), .Z(n1097) );
  CENXL U1446 ( .A(n1898), .B(n109), .Z(n1096) );
  CENXL U1447 ( .A(n109), .B(n1407), .Z(n1094) );
  CENXL U1448 ( .A(n109), .B(n1408), .Z(n1095) );
  CENXL U1449 ( .A(n109), .B(a[30]), .Z(n114) );
  CANR1XL U1450 ( .A(n265), .B(n246), .C(n247), .Z(n1571) );
  CND2X1 U1451 ( .A(n1589), .B(n1581), .Z(n1574) );
  CND2X2 U1452 ( .A(n1572), .B(n1573), .Z(n1575) );
  CND2X2 U1453 ( .A(n1574), .B(n1575), .Z(n542) );
  CIVX2 U1454 ( .A(n1589), .Z(n1572) );
  CIVX2 U1455 ( .A(n1581), .Z(n1573) );
  COND2X2 U1456 ( .A(n36), .B(n1261), .C(n1260), .D(n1606), .Z(n977) );
  CEOX2 U1457 ( .A(n876), .B(n930), .Z(n1576) );
  CEOXL U1458 ( .A(n1576), .B(n1030), .Z(n404) );
  CND2XL U1459 ( .A(n1580), .B(n930), .Z(n1577) );
  CND2XL U1460 ( .A(n1580), .B(n876), .Z(n1578) );
  CND2XL U1461 ( .A(n930), .B(n876), .Z(n1579) );
  CND3XL U1462 ( .A(n1577), .B(n1578), .C(n1579), .Z(n403) );
  COND2XL U1463 ( .A(n18), .B(n1316), .C(n15), .D(n1315), .Z(n1580) );
  COND2XL U1464 ( .A(n18), .B(n1316), .C(n15), .D(n1315), .Z(n1030) );
  CND2X1 U1465 ( .A(n720), .B(n731), .Z(n276) );
  CND2X1 U1466 ( .A(n169), .B(n181), .Z(n167) );
  CNR2XL U1467 ( .A(n744), .B(n753), .Z(n1582) );
  CFA1X1 U1468 ( .A(n897), .B(n1007), .CI(n981), .CO(n531), .S(n532) );
  COND1X1 U1469 ( .A(n248), .B(n252), .C(n249), .Z(n247) );
  CNR2X2 U1470 ( .A(n720), .B(n731), .Z(n275) );
  COND1X1 U1471 ( .A(n176), .B(n184), .C(n179), .Z(n175) );
  CND2X2 U1472 ( .A(n567), .B(n1583), .Z(n1584) );
  CND2X2 U1473 ( .A(n1584), .B(n1585), .Z(n1589) );
  CIVX2 U1474 ( .A(n565), .Z(n1583) );
  CENXL U1475 ( .A(n1898), .B(n113), .Z(n1091) );
  CENXL U1476 ( .A(n113), .B(n1408), .Z(n1090) );
  CND2IXL U1477 ( .B(n1899), .A(n113), .Z(n1092) );
  CNR2X2 U1478 ( .A(n187), .B(n192), .Z(n181) );
  CIVXL U1479 ( .A(n1556), .Z(n217) );
  COND1XL U1480 ( .A(n214), .B(n231), .C(n1556), .Z(n213) );
  CFA1X1 U1481 ( .A(n879), .B(n1005), .CI(n933), .CO(n483), .S(n484) );
  CIVX1 U1482 ( .A(n256), .Z(n254) );
  CND3X1 U1483 ( .A(n1827), .B(n1828), .C(n1829), .Z(n563) );
  CNR2X1 U1484 ( .A(n604), .B(n623), .Z(n225) );
  CND2X4 U1485 ( .A(n1422), .B(n1606), .Z(n36) );
  COND2X1 U1486 ( .A(n36), .B(n1282), .C(n1281), .D(n1606), .Z(n998) );
  COND2X1 U1487 ( .A(n36), .B(n1280), .C(n1279), .D(n1606), .Z(n996) );
  COND2X2 U1488 ( .A(n36), .B(n1265), .C(n1264), .D(n1606), .Z(n981) );
  CEO3X1 U1489 ( .A(n1639), .B(n1722), .C(n1807), .Z(n552) );
  CND2X1 U1490 ( .A(n1639), .B(n1807), .Z(n1586) );
  CND2X1 U1491 ( .A(n1639), .B(n1722), .Z(n1587) );
  CND2X1 U1492 ( .A(n1807), .B(n1722), .Z(n1588) );
  CND3XL U1493 ( .A(n1586), .B(n1587), .C(n1588), .Z(n551) );
  CEO3X2 U1494 ( .A(n1735), .B(n552), .C(n571), .Z(n546) );
  CND2X1 U1495 ( .A(n1735), .B(n552), .Z(n1590) );
  CND3X2 U1496 ( .A(n1590), .B(n1591), .C(n1592), .Z(n545) );
  CND2XL U1497 ( .A(n567), .B(n565), .Z(n1593) );
  CND2X1 U1498 ( .A(n567), .B(n546), .Z(n1594) );
  CND2XL U1499 ( .A(n565), .B(n546), .Z(n1595) );
  CND3X1 U1500 ( .A(n1593), .B(n1594), .C(n1595), .Z(n541) );
  CND2X1 U1501 ( .A(n492), .B(n515), .Z(n188) );
  COND1X1 U1502 ( .A(n171), .B(n179), .C(n172), .Z(n170) );
  COND1XL U1503 ( .A(n251), .B(n264), .C(n252), .Z(n250) );
  COND2X1 U1504 ( .A(n53), .B(n1215), .C(n1214), .D(n50), .Z(n933) );
  CENXL U1505 ( .A(n1873), .B(n1392), .Z(n1214) );
  CND2X2 U1506 ( .A(n516), .B(n539), .Z(n193) );
  CIVXL U1507 ( .A(n176), .Z(n341) );
  CNR2X2 U1508 ( .A(n466), .B(n491), .Z(n176) );
  CND2X1 U1509 ( .A(n1638), .B(n1805), .Z(n1596) );
  CND2X1 U1510 ( .A(n1638), .B(n1700), .Z(n1597) );
  CND2X1 U1511 ( .A(n1805), .B(n1700), .Z(n1598) );
  CND3X2 U1512 ( .A(n1596), .B(n1597), .C(n1598), .Z(n613) );
  CANR1X1 U1513 ( .A(n196), .B(n232), .C(n197), .Z(n1599) );
  CANR1X1 U1514 ( .A(n196), .B(n232), .C(n197), .Z(n195) );
  CENXL U1515 ( .A(n224), .B(n128), .Z(product[22]) );
  CENXL U1516 ( .A(n204), .B(n126), .Z(product[24]) );
  COND1X1 U1517 ( .A(n305), .B(n293), .C(n294), .Z(n292) );
  CIVXL U1518 ( .A(n1286), .Z(n1601) );
  CIVXL U1519 ( .A(n1601), .Z(n1602) );
  CENXL U1520 ( .A(n1858), .B(b[26]), .Z(n1286) );
  CENXL U1521 ( .A(n194), .B(n125), .Z(product[25]) );
  CENXL U1522 ( .A(n1603), .B(n122), .Z(product[28]) );
  CAOR1X1 U1523 ( .A(n174), .B(n1548), .C(n175), .Z(n1603) );
  CENXL U1524 ( .A(n1604), .B(n189), .Z(product[26]) );
  CAN2XL U1525 ( .A(n342), .B(n188), .Z(n1604) );
  CNR2X2 U1526 ( .A(n492), .B(n515), .Z(n187) );
  COND2X1 U1527 ( .A(n53), .B(n1214), .C(n1213), .D(n50), .Z(n932) );
  CNR2X2 U1528 ( .A(n516), .B(n539), .Z(n192) );
  CANR1X2 U1529 ( .A(n284), .B(n292), .C(n285), .Z(n283) );
  CIVXL U1530 ( .A(n232), .Z(n231) );
  CFA1XL U1531 ( .A(n848), .B(n870), .CI(n858), .CO(n601), .S(n602) );
  CENXL U1532 ( .A(n1869), .B(n1386), .Z(n1233) );
  COND2X2 U1533 ( .A(n36), .B(n1262), .C(n1261), .D(n1606), .Z(n978) );
  COND1X1 U1534 ( .A(n233), .B(n245), .C(n234), .Z(n232) );
  CIVXL U1535 ( .A(n1571), .Z(n244) );
  COND2X2 U1536 ( .A(n44), .B(n1235), .C(n1234), .D(n1836), .Z(n952) );
  CFA1XL U1537 ( .A(n847), .B(n883), .CI(n869), .CO(n579), .S(n580) );
  CFA1XL U1538 ( .A(n860), .B(n886), .CI(n872), .CO(n639), .S(n640) );
  CENXL U1539 ( .A(n166), .B(n121), .Z(product[29]) );
  CANR1X1 U1540 ( .A(n1609), .B(n166), .C(n1610), .Z(n152) );
  CANR1X1 U1541 ( .A(n1614), .B(n166), .C(n163), .Z(n161) );
  COND2XL U1542 ( .A(n44), .B(n1241), .C(n1240), .D(n1836), .Z(n958) );
  CIVX1 U1543 ( .A(n1599), .Z(n194) );
  CANR1X1 U1544 ( .A(n246), .B(n265), .C(n247), .Z(n245) );
  COND1X1 U1545 ( .A(n283), .B(n266), .C(n267), .Z(n265) );
  COND1X1 U1546 ( .A(n311), .B(n313), .C(n312), .Z(n310) );
  CANR1X1 U1547 ( .A(n318), .B(n1628), .C(n315), .Z(n313) );
  CND2IX1 U1548 ( .B(n1608), .A(n74), .Z(n77) );
  CENX1 U1549 ( .A(a[16]), .B(n1883), .Z(n1608) );
  CENX1 U1550 ( .A(n1876), .B(n1393), .Z(n1192) );
  CENX1 U1551 ( .A(n1864), .B(n1393), .Z(n1267) );
  CENX1 U1552 ( .A(n1880), .B(n1393), .Z(n1171) );
  CENX1 U1553 ( .A(n1850), .B(n1393), .Z(n1327) );
  CENX1 U1554 ( .A(n142), .B(n310), .Z(product[8]) );
  CNIVX1 U1555 ( .A(n1397), .Z(n1846) );
  COND2XL U1556 ( .A(n69), .B(n1175), .C(n1174), .D(n66), .Z(n895) );
  CNR2IXL U1557 ( .B(n1899), .A(n58), .Z(n928) );
  CND2IX4 U1558 ( .B(n1607), .A(n66), .Z(n69) );
  CENXL U1559 ( .A(a[14]), .B(n1879), .Z(n1607) );
  CND2X2 U1560 ( .A(n1423), .B(n24), .Z(n27) );
  CNIVX1 U1561 ( .A(n42), .Z(n1836) );
  CENX1 U1562 ( .A(n146), .B(n326), .Z(product[4]) );
  CND2XL U1563 ( .A(n1614), .B(n165), .Z(n121) );
  CNR2IXL U1564 ( .B(n181), .A(n176), .Z(n174) );
  CND2XL U1565 ( .A(n1618), .B(n1619), .Z(n233) );
  CND2XL U1566 ( .A(n273), .B(n1620), .Z(n266) );
  CIVX1 U1567 ( .A(n223), .Z(n221) );
  CEOXL U1568 ( .A(n130), .B(n239), .Z(product[20]) );
  CND2XL U1569 ( .A(n1618), .B(n238), .Z(n130) );
  CEOXL U1570 ( .A(n136), .B(n277), .Z(product[14]) );
  CEOXL U1571 ( .A(n135), .B(n272), .Z(product[15]) );
  CND2XL U1572 ( .A(n1620), .B(n271), .Z(n135) );
  CNR2XL U1573 ( .A(n275), .B(n280), .Z(n273) );
  CEOXL U1574 ( .A(n134), .B(n264), .Z(product[16]) );
  CND2XL U1575 ( .A(n352), .B(n259), .Z(n134) );
  CND2XL U1576 ( .A(n216), .B(n1611), .Z(n205) );
  CND2XL U1577 ( .A(n1619), .B(n243), .Z(n131) );
  CND2XL U1578 ( .A(n355), .B(n281), .Z(n137) );
  CND2XL U1579 ( .A(n1617), .B(n352), .Z(n251) );
  COR2XL U1580 ( .A(n412), .B(n439), .Z(n1614) );
  CNR2XL U1581 ( .A(n286), .B(n289), .Z(n284) );
  CND2XL U1582 ( .A(n383), .B(n368), .Z(n151) );
  CND2XL U1583 ( .A(n744), .B(n753), .Z(n287) );
  CNIVX2 U1584 ( .A(n1396), .Z(n1847) );
  CND2IXL U1585 ( .B(n311), .A(n312), .Z(n143) );
  CND2XL U1586 ( .A(n1626), .B(n298), .Z(n140) );
  CND2XL U1587 ( .A(n357), .B(n290), .Z(n139) );
  CND2XL U1588 ( .A(n1627), .B(n309), .Z(n142) );
  CND2XL U1589 ( .A(n1625), .B(n303), .Z(n141) );
  CND2XL U1590 ( .A(n356), .B(n287), .Z(n138) );
  CNR2XL U1591 ( .A(n796), .B(n799), .Z(n319) );
  CND2XL U1592 ( .A(n585), .B(n564), .Z(n1832) );
  CND2XL U1593 ( .A(n800), .B(n801), .Z(n325) );
  CNR2IXL U1594 ( .B(n1899), .A(n82), .Z(n874) );
  COND2XL U1595 ( .A(n84), .B(n1148), .C(n1147), .D(n82), .Z(n870) );
  CIVX2 U1596 ( .A(n1866), .Z(n1863) );
  CND2X4 U1597 ( .A(n1424), .B(n15), .Z(n18) );
  CIVX1 U1598 ( .A(n1874), .Z(n1873) );
  COND2XL U1599 ( .A(n36), .B(n1279), .C(n1278), .D(n1606), .Z(n995) );
  COND2XL U1600 ( .A(n44), .B(n1254), .C(n1253), .D(n1836), .Z(n971) );
  COND2XL U1601 ( .A(n44), .B(n1247), .C(n1246), .D(n1836), .Z(n964) );
  COND2XL U1602 ( .A(n44), .B(n1244), .C(n1243), .D(n1836), .Z(n961) );
  COR2XL U1603 ( .A(n772), .B(n779), .Z(n1625) );
  COND2XL U1604 ( .A(n18), .B(n1342), .C(n15), .D(n1341), .Z(n1056) );
  COND2XL U1605 ( .A(n18), .B(n1343), .C(n15), .D(n1342), .Z(n1057) );
  COND2XL U1606 ( .A(n27), .B(n1312), .C(n24), .D(n1311), .Z(n1027) );
  COND2XL U1607 ( .A(n84), .B(n1143), .C(n1142), .D(n82), .Z(n865) );
  COND2XL U1608 ( .A(n53), .B(n1230), .C(n1229), .D(n50), .Z(n948) );
  COND2XL U1609 ( .A(n84), .B(n1150), .C(n1149), .D(n82), .Z(n872) );
  COND2XL U1610 ( .A(n84), .B(n1147), .C(n1146), .D(n82), .Z(n869) );
  COND2XL U1611 ( .A(n53), .B(n1228), .C(n1227), .D(n50), .Z(n946) );
  COND2XL U1612 ( .A(n18), .B(n1340), .C(n15), .D(n1339), .Z(n1054) );
  COND2XL U1613 ( .A(n84), .B(n1151), .C(n1150), .D(n82), .Z(n873) );
  COND2XL U1614 ( .A(n84), .B(n1149), .C(n1148), .D(n82), .Z(n871) );
  CND2XL U1615 ( .A(n1628), .B(n317), .Z(n144) );
  CNR2IXL U1616 ( .B(n1899), .A(n6), .Z(product[0]) );
  COND1X1 U1617 ( .A(n1816), .B(n1818), .C(n1817), .Z(n326) );
  COND1X1 U1618 ( .A(n321), .B(n1821), .C(n1820), .Z(n318) );
  CEOXL U1619 ( .A(a[8]), .B(n1870), .Z(n1421) );
  CENX1 U1620 ( .A(n1872), .B(a[12]), .Z(n58) );
  CENX1 U1621 ( .A(n1875), .B(a[14]), .Z(n66) );
  CEOXL U1622 ( .A(a[12]), .B(n1876), .Z(n1605) );
  CND2X1 U1623 ( .A(n89), .B(n1415), .Z(n91) );
  COND2XL U1624 ( .A(n102), .B(n1110), .C(n1109), .D(n100), .Z(n835) );
  CIVXL U1625 ( .A(n104), .Z(n1437) );
  CEOXL U1626 ( .A(a[30]), .B(a[31]), .Z(n1410) );
  CIVXL U1627 ( .A(n99), .Z(n1897) );
  CND2IXL U1628 ( .B(n1821), .A(n1820), .Z(n145) );
  CND2XL U1629 ( .A(n1822), .B(n1819), .Z(n146) );
  CANR1XL U1630 ( .A(n1611), .B(n217), .C(n210), .Z(n206) );
  CND2X1 U1631 ( .A(n1611), .B(n212), .Z(n127) );
  CND2X1 U1632 ( .A(n1551), .B(n347), .Z(n214) );
  CAOR1X1 U1633 ( .A(n163), .B(n1613), .C(n158), .Z(n1610) );
  CENX1 U1634 ( .A(n1867), .B(n1389), .Z(n1236) );
  CENX1 U1635 ( .A(n1867), .B(n1553), .Z(n1237) );
  CENX1 U1636 ( .A(n1868), .B(n1550), .Z(n1238) );
  CENX1 U1637 ( .A(n1867), .B(n1387), .Z(n1234) );
  CENX1 U1638 ( .A(n1870), .B(n1848), .Z(n1242) );
  CENX1 U1639 ( .A(n1868), .B(n1849), .Z(n1241) );
  CENX1 U1640 ( .A(n1870), .B(n1845), .Z(n1245) );
  CENX1 U1641 ( .A(n1867), .B(n1847), .Z(n1243) );
  CNR2X1 U1642 ( .A(n440), .B(n465), .Z(n171) );
  CENX1 U1643 ( .A(n257), .B(n133), .Z(product[17]) );
  CND2X1 U1644 ( .A(n1617), .B(n256), .Z(n133) );
  COND1XL U1645 ( .A(n258), .B(n264), .C(n259), .Z(n257) );
  CENX1 U1646 ( .A(n250), .B(n132), .Z(product[18]) );
  CND2X1 U1647 ( .A(n350), .B(n249), .Z(n132) );
  CENX1 U1648 ( .A(n244), .B(n131), .Z(product[19]) );
  COND1XL U1649 ( .A(n225), .B(n231), .C(n226), .Z(n224) );
  CENX1 U1650 ( .A(n282), .B(n137), .Z(product[13]) );
  COND1XL U1651 ( .A(n205), .B(n231), .C(n206), .Z(n204) );
  COR2X1 U1652 ( .A(n562), .B(n583), .Z(n1611) );
  CND2X1 U1653 ( .A(n354), .B(n276), .Z(n136) );
  CANR1XL U1654 ( .A(n355), .B(n282), .C(n279), .Z(n277) );
  CANR1XL U1655 ( .A(n273), .B(n282), .C(n274), .Z(n272) );
  CANR1XL U1656 ( .A(n1619), .B(n244), .C(n241), .Z(n239) );
  CEOXL U1657 ( .A(n129), .B(n231), .Z(product[21]) );
  CND2XL U1658 ( .A(n347), .B(n226), .Z(n129) );
  COR2X1 U1659 ( .A(n584), .B(n603), .Z(n1612) );
  COR2X1 U1660 ( .A(n384), .B(n411), .Z(n1613) );
  CND2X1 U1661 ( .A(n562), .B(n583), .Z(n212) );
  CND2X1 U1662 ( .A(n584), .B(n603), .Z(n223) );
  CND2X1 U1663 ( .A(n412), .B(n439), .Z(n165) );
  CND2X1 U1664 ( .A(n384), .B(n411), .Z(n160) );
  CND2X1 U1665 ( .A(n466), .B(n491), .Z(n179) );
  CENX1 U1666 ( .A(n1861), .B(n1386), .Z(n1260) );
  CENX1 U1667 ( .A(n1851), .B(n1386), .Z(n1320) );
  CENX1 U1668 ( .A(n1855), .B(n1386), .Z(n1289) );
  CENX1 U1669 ( .A(n1861), .B(n1554), .Z(n1264) );
  CENX1 U1670 ( .A(n1861), .B(n1387), .Z(n1261) );
  CENX1 U1671 ( .A(n1862), .B(n1389), .Z(n1263) );
  CENX1 U1672 ( .A(n1872), .B(n1389), .Z(n1211) );
  CENX1 U1673 ( .A(n1872), .B(n1555), .Z(n1212) );
  CENX1 U1674 ( .A(n1876), .B(n1392), .Z(n1191) );
  CENX1 U1675 ( .A(n1864), .B(n1392), .Z(n1266) );
  CENX1 U1676 ( .A(n1855), .B(n1389), .Z(n1292) );
  CENX1 U1677 ( .A(n1850), .B(n1555), .Z(n1324) );
  CENX1 U1678 ( .A(n1858), .B(n1555), .Z(n1293) );
  CENX1 U1679 ( .A(n1615), .B(n564), .Z(n562) );
  CENX1 U1680 ( .A(n566), .B(n585), .Z(n1615) );
  CENX1 U1681 ( .A(n288), .B(n138), .Z(product[12]) );
  COND1XL U1682 ( .A(n289), .B(n291), .C(n290), .Z(n288) );
  CENX1 U1683 ( .A(n1863), .B(b[25]), .Z(n1258) );
  CENX1 U1684 ( .A(n1876), .B(n1555), .Z(n1189) );
  CENX1 U1685 ( .A(n1880), .B(n1392), .Z(n1170) );
  CENX1 U1686 ( .A(n1864), .B(n1848), .Z(n1269) );
  CENX1 U1687 ( .A(n1862), .B(n1550), .Z(n1265) );
  CENX1 U1688 ( .A(n1873), .B(n1849), .Z(n1216) );
  CENX1 U1689 ( .A(n1880), .B(n1846), .Z(n1175) );
  CENX1 U1690 ( .A(n1864), .B(n1847), .Z(n1270) );
  CENX1 U1691 ( .A(n1873), .B(n1846), .Z(n1219) );
  CENX1 U1692 ( .A(n1864), .B(n1849), .Z(n1268) );
  CENX1 U1693 ( .A(n1880), .B(n1847), .Z(n1174) );
  CENX1 U1694 ( .A(n1872), .B(n1847), .Z(n1218) );
  CENX1 U1695 ( .A(n1888), .B(n1843), .Z(n1142) );
  CNR2X1 U1696 ( .A(n744), .B(n753), .Z(n286) );
  CENX1 U1697 ( .A(n1616), .B(n442), .Z(n440) );
  CENX1 U1698 ( .A(n444), .B(n467), .Z(n1616) );
  CENX1 U1699 ( .A(n1876), .B(n1550), .Z(n1190) );
  CENX1 U1700 ( .A(n1880), .B(n1843), .Z(n1178) );
  CENX1 U1701 ( .A(n1875), .B(n1845), .Z(n1197) );
  CENX1 U1702 ( .A(n1873), .B(n1848), .Z(n1217) );
  CENX1 U1703 ( .A(n1880), .B(n1844), .Z(n1177) );
  CENX1 U1704 ( .A(n1880), .B(n1845), .Z(n1176) );
  CENX1 U1705 ( .A(n1876), .B(n1848), .Z(n1194) );
  CENX1 U1706 ( .A(n1876), .B(n1849), .Z(n1193) );
  CENX1 U1707 ( .A(n1879), .B(n1848), .Z(n1173) );
  CENX1 U1708 ( .A(n1879), .B(n1849), .Z(n1172) );
  CENX1 U1709 ( .A(n1884), .B(n1848), .Z(n1154) );
  CENX1 U1710 ( .A(n1862), .B(n1843), .Z(n1274) );
  CENX1 U1711 ( .A(n1862), .B(n1844), .Z(n1273) );
  CENX1 U1712 ( .A(n1864), .B(n1845), .Z(n1272) );
  CENX1 U1713 ( .A(n1864), .B(n1846), .Z(n1271) );
  CENX1 U1714 ( .A(n1873), .B(n1843), .Z(n1222) );
  CENX1 U1715 ( .A(n1873), .B(n1844), .Z(n1221) );
  CENX1 U1716 ( .A(n1873), .B(n1845), .Z(n1220) );
  CENX1 U1717 ( .A(n1876), .B(n1846), .Z(n1196) );
  CENX1 U1718 ( .A(n1876), .B(n1847), .Z(n1195) );
  CENX1 U1719 ( .A(n1884), .B(n1843), .Z(n1159) );
  CENX1 U1720 ( .A(n1884), .B(n1844), .Z(n1158) );
  CENX1 U1721 ( .A(n1884), .B(n1845), .Z(n1157) );
  CENX1 U1722 ( .A(n1888), .B(n1844), .Z(n1141) );
  CENX1 U1723 ( .A(n1884), .B(n1846), .Z(n1156) );
  CENX1 U1724 ( .A(n1892), .B(n1843), .Z(n1127) );
  CENX1 U1725 ( .A(n1888), .B(n1845), .Z(n1140) );
  CENX1 U1726 ( .A(n1884), .B(n1847), .Z(n1155) );
  CENX1 U1727 ( .A(n1892), .B(n1844), .Z(n1126) );
  CENX1 U1728 ( .A(n1887), .B(n1846), .Z(n1139) );
  CENX1 U1729 ( .A(n1869), .B(n1844), .Z(n1246) );
  CENX1 U1730 ( .A(n1870), .B(n1843), .Z(n1247) );
  CENX1 U1731 ( .A(n1870), .B(n1846), .Z(n1244) );
  CENX1 U1732 ( .A(n1850), .B(b[26]), .Z(n1317) );
  CENX1 U1733 ( .A(n1851), .B(n1550), .Z(n1325) );
  CENX1 U1734 ( .A(n1859), .B(n1550), .Z(n1294) );
  CENX1 U1735 ( .A(n1853), .B(n1848), .Z(n1329) );
  CENX1 U1736 ( .A(n1853), .B(n1849), .Z(n1328) );
  CENX1 U1737 ( .A(n1855), .B(n1848), .Z(n1298) );
  CENX1 U1738 ( .A(n1850), .B(n1843), .Z(n1334) );
  CENX1 U1739 ( .A(n1853), .B(n1846), .Z(n1331) );
  CENX1 U1740 ( .A(n1853), .B(n1847), .Z(n1330) );
  CENX1 U1741 ( .A(n1851), .B(n1387), .Z(n1321) );
  CENX1 U1742 ( .A(n1855), .B(n1387), .Z(n1290) );
  CENX1 U1743 ( .A(n1853), .B(b[24]), .Z(n1319) );
  CENX1 U1744 ( .A(n1858), .B(b[24]), .Z(n1288) );
  CENX1 U1745 ( .A(n1850), .B(b[25]), .Z(n1318) );
  CENX1 U1746 ( .A(n1858), .B(b[25]), .Z(n1287) );
  CENX1 U1747 ( .A(n1853), .B(n1844), .Z(n1333) );
  CENX1 U1748 ( .A(n1851), .B(n1845), .Z(n1332) );
  CENX1 U1749 ( .A(n1857), .B(n1843), .Z(n1303) );
  CENX1 U1750 ( .A(n1858), .B(n1844), .Z(n1302) );
  CENX1 U1751 ( .A(n1858), .B(n1845), .Z(n1301) );
  CENX1 U1752 ( .A(n1858), .B(n1846), .Z(n1300) );
  CENX1 U1753 ( .A(n1858), .B(n1847), .Z(n1299) );
  CENX1 U1754 ( .A(n1855), .B(n1849), .Z(n1297) );
  CNR2X1 U1755 ( .A(n732), .B(n743), .Z(n280) );
  CENX1 U1756 ( .A(n1873), .B(n1550), .Z(n1213) );
  CENX1 U1757 ( .A(n1884), .B(n1849), .Z(n1153) );
  CENX1 U1758 ( .A(n1894), .B(n1843), .Z(n1114) );
  CENX1 U1759 ( .A(n1892), .B(n1845), .Z(n1125) );
  CENX1 U1760 ( .A(n1887), .B(n1847), .Z(n1138) );
  CENX1 U1761 ( .A(n1852), .B(b[29]), .Z(n1314) );
  CENX1 U1762 ( .A(n141), .B(n304), .Z(product[9]) );
  CND3XL U1763 ( .A(n1830), .B(n1831), .C(n1832), .Z(n561) );
  CNR2X1 U1764 ( .A(n692), .B(n705), .Z(n258) );
  CEOX1 U1765 ( .A(n299), .B(n140), .Z(product[10]) );
  CANR1XL U1766 ( .A(n1625), .B(n304), .C(n301), .Z(n299) );
  CEOX1 U1767 ( .A(n139), .B(n291), .Z(product[11]) );
  COR2X1 U1768 ( .A(n676), .B(n691), .Z(n1617) );
  COR2X1 U1769 ( .A(n624), .B(n641), .Z(n1618) );
  COR2X1 U1770 ( .A(n642), .B(n659), .Z(n1619) );
  COR2X1 U1771 ( .A(n706), .B(n719), .Z(n1620) );
  CND2X1 U1772 ( .A(n692), .B(n705), .Z(n259) );
  CND2X1 U1773 ( .A(n732), .B(n743), .Z(n281) );
  CND2X1 U1774 ( .A(n604), .B(n623), .Z(n226) );
  CNIVX1 U1775 ( .A(n1398), .Z(n1845) );
  CND2X1 U1776 ( .A(n642), .B(n659), .Z(n243) );
  CND2X1 U1777 ( .A(n676), .B(n691), .Z(n256) );
  CND2X1 U1778 ( .A(n706), .B(n719), .Z(n271) );
  CND2X1 U1779 ( .A(n624), .B(n641), .Z(n238) );
  CND2X1 U1780 ( .A(n1088), .B(n1058), .Z(n333) );
  CNR2X1 U1781 ( .A(n802), .B(n817), .Z(n327) );
  CNIVX1 U1782 ( .A(n1394), .Z(n1849) );
  CND2X1 U1783 ( .A(n660), .B(n675), .Z(n249) );
  COR2X1 U1784 ( .A(n540), .B(n561), .Z(n1621) );
  COR2X1 U1785 ( .A(n1088), .B(n1058), .Z(n1622) );
  CND2X1 U1786 ( .A(n540), .B(n561), .Z(n203) );
  COR2X1 U1787 ( .A(n383), .B(n368), .Z(n1623) );
  CND2XL U1788 ( .A(n796), .B(n799), .Z(n320) );
  CND2X1 U1789 ( .A(n802), .B(n817), .Z(n328) );
  COR2X1 U1790 ( .A(n800), .B(n801), .Z(n1624) );
  CIVX2 U1791 ( .A(n1877), .Z(n1875) );
  CENX1 U1792 ( .A(n1868), .B(n1838), .Z(n1252) );
  CENX1 U1793 ( .A(n1850), .B(n1838), .Z(n1339) );
  CENX1 U1794 ( .A(n1856), .B(n1838), .Z(n1308) );
  CIVX2 U1795 ( .A(n1895), .Z(n1894) );
  CNR2IX1 U1796 ( .B(n1899), .A(n66), .Z(n908) );
  CNR2IX1 U1797 ( .B(n1899), .A(n1606), .Z(n1000) );
  CNR2IXL U1798 ( .B(n1899), .A(n50), .Z(n950) );
  CNR2IX1 U1799 ( .B(n1899), .A(n114), .Z(n820) );
  COND2X1 U1800 ( .A(n107), .B(n1100), .C(n1099), .D(n105), .Z(n826) );
  CIVX2 U1801 ( .A(n1897), .Z(n1896) );
  CEOX1 U1802 ( .A(a[2]), .B(n1851), .Z(n1424) );
  CENX1 U1803 ( .A(n1863), .B(n1898), .Z(n1283) );
  CENX1 U1804 ( .A(n1868), .B(n1898), .Z(n1256) );
  CENX1 U1805 ( .A(n1872), .B(n1898), .Z(n1231) );
  CENX1 U1806 ( .A(n1879), .B(n1898), .Z(n1187) );
  CENX1 U1807 ( .A(n1898), .B(n1884), .Z(n1168) );
  CENX1 U1808 ( .A(n1898), .B(n1892), .Z(n1136) );
  CENX1 U1809 ( .A(n1883), .B(n1837), .Z(n1165) );
  CENX1 U1810 ( .A(n1882), .B(n1840), .Z(n1162) );
  CENX1 U1811 ( .A(n1894), .B(n1837), .Z(n1120) );
  CENX1 U1812 ( .A(n1894), .B(n1838), .Z(n1119) );
  CENX1 U1813 ( .A(n1896), .B(n1838), .Z(n1108) );
  CENX1 U1814 ( .A(n1887), .B(n1837), .Z(n1148) );
  CENX1 U1815 ( .A(n1896), .B(n1837), .Z(n1109) );
  CIVX1 U1816 ( .A(n1877), .Z(n1876) );
  CENX1 U1817 ( .A(n1898), .B(n1896), .Z(n1112) );
  CENX1 U1818 ( .A(n1875), .B(n1840), .Z(n1202) );
  CENX1 U1819 ( .A(n1880), .B(n1841), .Z(n1180) );
  CENX1 U1820 ( .A(n1878), .B(n1839), .Z(n1182) );
  CENX1 U1821 ( .A(n1882), .B(n1839), .Z(n1163) );
  CENX1 U1822 ( .A(n1890), .B(n1840), .Z(n1130) );
  CENX1 U1823 ( .A(n1888), .B(n1842), .Z(n1143) );
  CENX1 U1824 ( .A(n1891), .B(n1837), .Z(n1133) );
  COND2XL U1825 ( .A(n91), .B(n1893), .C(n1137), .D(n89), .Z(n808) );
  CENX1 U1826 ( .A(n1878), .B(n1840), .Z(n1181) );
  CENX1 U1827 ( .A(n1880), .B(n1842), .Z(n1179) );
  CENX1 U1828 ( .A(n1886), .B(n1839), .Z(n1146) );
  CENX1 U1829 ( .A(n1875), .B(n1842), .Z(n1200) );
  CENX1 U1830 ( .A(n1884), .B(n1841), .Z(n1161) );
  CENX1 U1831 ( .A(n1891), .B(n1841), .Z(n1129) );
  CENX1 U1832 ( .A(n1894), .B(n1839), .Z(n1118) );
  CENX1 U1833 ( .A(n1862), .B(n1839), .Z(n1278) );
  CNR2X1 U1834 ( .A(n754), .B(n763), .Z(n289) );
  CNR2IX1 U1835 ( .B(n1899), .A(n15), .Z(n1058) );
  CENX1 U1836 ( .A(n1875), .B(n1841), .Z(n1201) );
  CENX1 U1837 ( .A(n1886), .B(n1838), .Z(n1147) );
  CENX1 U1838 ( .A(n1898), .B(n1894), .Z(n1123) );
  CENX1 U1839 ( .A(n1875), .B(n1837), .Z(n1205) );
  CENX1 U1840 ( .A(n1875), .B(n1839), .Z(n1203) );
  CENX1 U1841 ( .A(n1872), .B(n1837), .Z(n1228) );
  CENX1 U1842 ( .A(n1868), .B(n1839), .Z(n1251) );
  CENX1 U1843 ( .A(n1862), .B(n1841), .Z(n1276) );
  CENX1 U1844 ( .A(n1864), .B(n1842), .Z(n1275) );
  CENX1 U1845 ( .A(n1868), .B(n1840), .Z(n1250) );
  CENX1 U1846 ( .A(n1868), .B(n1841), .Z(n1249) );
  CENX1 U1847 ( .A(n1872), .B(n1840), .Z(n1225) );
  CENX1 U1848 ( .A(n1879), .B(n1837), .Z(n1184) );
  CENX1 U1849 ( .A(n1872), .B(n1841), .Z(n1224) );
  CENX1 U1850 ( .A(n1873), .B(n1842), .Z(n1223) );
  CENX1 U1851 ( .A(n1886), .B(n1840), .Z(n1145) );
  CENX1 U1852 ( .A(n1883), .B(n1842), .Z(n1160) );
  CENX1 U1853 ( .A(n1890), .B(n1839), .Z(n1131) );
  CENX1 U1854 ( .A(n1887), .B(n1841), .Z(n1144) );
  CENX1 U1855 ( .A(n1894), .B(n1840), .Z(n1117) );
  CENX1 U1856 ( .A(n1892), .B(n1842), .Z(n1128) );
  CENX1 U1857 ( .A(n1894), .B(n1841), .Z(n1116) );
  CENX1 U1858 ( .A(n1896), .B(n1840), .Z(n1106) );
  CENX1 U1859 ( .A(n1869), .B(n1842), .Z(n1248) );
  CENX1 U1860 ( .A(n1894), .B(n1842), .Z(n1115) );
  CENX1 U1861 ( .A(n1867), .B(n1837), .Z(n1253) );
  CENX1 U1862 ( .A(n1872), .B(n1839), .Z(n1226) );
  CENX1 U1863 ( .A(n1850), .B(n1837), .Z(n1340) );
  CENX1 U1864 ( .A(n1851), .B(n1839), .Z(n1338) );
  CENX1 U1865 ( .A(n1851), .B(n1840), .Z(n1337) );
  CENX1 U1866 ( .A(n1851), .B(n1841), .Z(n1336) );
  CENX1 U1867 ( .A(n1851), .B(n1842), .Z(n1335) );
  CENX1 U1868 ( .A(n1858), .B(n1837), .Z(n1309) );
  CENX1 U1869 ( .A(n1856), .B(n1839), .Z(n1307) );
  CENX1 U1870 ( .A(n1856), .B(n1840), .Z(n1306) );
  CENX1 U1871 ( .A(n1856), .B(n1841), .Z(n1305) );
  CENX1 U1872 ( .A(n1857), .B(n1842), .Z(n1304) );
  CIVX2 U1873 ( .A(n1874), .Z(n1872) );
  CENX1 U1874 ( .A(n1896), .B(n1841), .Z(n1105) );
  CENX1 U1875 ( .A(n1875), .B(n1899), .Z(n1208) );
  CENX1 U1876 ( .A(n1857), .B(n1899), .Z(n1312) );
  CNR2IX1 U1877 ( .B(n1899), .A(n24), .Z(n1028) );
  CENX1 U1878 ( .A(n1852), .B(n1898), .Z(n1343) );
  CNR2X1 U1879 ( .A(n786), .B(n791), .Z(n311) );
  COR2X1 U1880 ( .A(n764), .B(n771), .Z(n1626) );
  CNR2IX1 U1881 ( .B(n1899), .A(n105), .Z(n830) );
  COND2X1 U1882 ( .A(n102), .B(n1111), .C(n1110), .D(n100), .Z(n836) );
  COND2X1 U1883 ( .A(n97), .B(n1120), .C(n1119), .D(n95), .Z(n844) );
  CNIVX1 U1884 ( .A(n1400), .Z(n1843) );
  COND2X1 U1885 ( .A(n107), .B(n1101), .C(n1100), .D(n105), .Z(n827) );
  COND2X1 U1886 ( .A(n102), .B(n1108), .C(n1107), .D(n100), .Z(n833) );
  CND2X1 U1887 ( .A(n754), .B(n763), .Z(n290) );
  CND2X1 U1888 ( .A(n772), .B(n779), .Z(n303) );
  CND2X1 U1889 ( .A(n780), .B(n785), .Z(n309) );
  CND2X1 U1890 ( .A(n764), .B(n771), .Z(n298) );
  CNIVX1 U1891 ( .A(n1399), .Z(n1844) );
  COR2X1 U1892 ( .A(n780), .B(n785), .Z(n1627) );
  CEOX1 U1893 ( .A(n825), .B(n831), .Z(n382) );
  COND2X1 U1894 ( .A(n107), .B(n1099), .C(n1098), .D(n105), .Z(n825) );
  CND2X1 U1895 ( .A(n786), .B(n791), .Z(n312) );
  CNR2IX1 U1896 ( .B(n1899), .A(n1836), .Z(n974) );
  COND2XL U1897 ( .A(n77), .B(n1163), .C(n1162), .D(n74), .Z(n884) );
  COND2XL U1898 ( .A(n53), .B(n1219), .C(n1218), .D(n50), .Z(n937) );
  COND2X1 U1899 ( .A(n36), .B(n1270), .C(n1269), .D(n1606), .Z(n986) );
  COND2XL U1900 ( .A(n69), .B(n1182), .C(n1181), .D(n66), .Z(n902) );
  COND2XL U1901 ( .A(n77), .B(n1167), .C(n1166), .D(n74), .Z(n888) );
  COND2XL U1902 ( .A(n77), .B(n1166), .C(n1165), .D(n74), .Z(n887) );
  CNR2IXL U1903 ( .B(n1899), .A(n89), .Z(n860) );
  COND2XL U1904 ( .A(n77), .B(n1165), .C(n1164), .D(n74), .Z(n886) );
  COND2X1 U1905 ( .A(n97), .B(n1123), .C(n1122), .D(n95), .Z(n847) );
  COND2XL U1906 ( .A(n77), .B(n1162), .C(n1161), .D(n74), .Z(n883) );
  CNR2IX1 U1907 ( .B(n1899), .A(n100), .Z(n838) );
  COND2X1 U1908 ( .A(n97), .B(n1122), .C(n1121), .D(n95), .Z(n846) );
  COND2XL U1909 ( .A(n91), .B(n1133), .C(n1132), .D(n89), .Z(n856) );
  COND2X1 U1910 ( .A(n1103), .B(n107), .C(n1102), .D(n105), .Z(n829) );
  COND2X1 U1911 ( .A(n97), .B(n1119), .C(n1118), .D(n95), .Z(n843) );
  COND2XL U1912 ( .A(n91), .B(n1130), .C(n1129), .D(n89), .Z(n853) );
  COND2X1 U1913 ( .A(n36), .B(n1269), .C(n1268), .D(n1606), .Z(n985) );
  CNR2IXL U1914 ( .B(n1899), .A(n74), .Z(n890) );
  COND2X1 U1915 ( .A(n61), .B(n1202), .C(n1201), .D(n58), .Z(n921) );
  COND2X1 U1916 ( .A(n69), .B(n1180), .C(n1179), .D(n66), .Z(n900) );
  COND2X1 U1917 ( .A(n61), .B(n1199), .C(n1198), .D(n58), .Z(n918) );
  CNR2IX1 U1918 ( .B(n1899), .A(n95), .Z(n848) );
  COND2XL U1919 ( .A(n91), .B(n1135), .C(n1134), .D(n89), .Z(n858) );
  COND2X1 U1920 ( .A(n97), .B(n1121), .C(n1120), .D(n95), .Z(n845) );
  CNR2IX1 U1921 ( .B(n1899), .A(n110), .Z(n824) );
  COND2X1 U1922 ( .A(n107), .B(n1102), .C(n1101), .D(n105), .Z(n828) );
  COND2X1 U1923 ( .A(n102), .B(n1109), .C(n1108), .D(n100), .Z(n834) );
  CENX1 U1924 ( .A(n144), .B(n318), .Z(product[6]) );
  CENX1 U1925 ( .A(n1882), .B(a[18]), .Z(n82) );
  CENX1 U1926 ( .A(n1890), .B(a[22]), .Z(n95) );
  CENX1 U1927 ( .A(n1894), .B(a[24]), .Z(n100) );
  CENX1 U1928 ( .A(n1896), .B(a[26]), .Z(n105) );
  CENX1 U1929 ( .A(n1875), .B(n1408), .Z(n1207) );
  CENX1 U1930 ( .A(n1863), .B(n1408), .Z(n1282) );
  CENX1 U1931 ( .A(n1868), .B(n1408), .Z(n1255) );
  CENX1 U1932 ( .A(n1872), .B(n1408), .Z(n1230) );
  CENX1 U1933 ( .A(n1872), .B(n1407), .Z(n1229) );
  CENX1 U1934 ( .A(n1862), .B(n1407), .Z(n1281) );
  CENX1 U1935 ( .A(n1867), .B(n1407), .Z(n1254) );
  CENX1 U1936 ( .A(n1852), .B(n1408), .Z(n1342) );
  CENX1 U1937 ( .A(n1853), .B(n1407), .Z(n1341) );
  CENX1 U1938 ( .A(n1855), .B(n1408), .Z(n1311) );
  CENX1 U1939 ( .A(n1856), .B(n1407), .Z(n1310) );
  CENX1 U1940 ( .A(n1887), .B(n1408), .Z(n1150) );
  CENX1 U1941 ( .A(n1894), .B(n1408), .Z(n1122) );
  CENX1 U1942 ( .A(n1887), .B(n1407), .Z(n1149) );
  CND2X1 U1943 ( .A(n100), .B(n1413), .Z(n102) );
  CEOXL U1944 ( .A(a[24]), .B(n1896), .Z(n1413) );
  CANR1XL U1945 ( .A(n326), .B(n1822), .C(n323), .Z(n321) );
  CND2X1 U1946 ( .A(n1412), .B(n105), .Z(n107) );
  CEOXL U1947 ( .A(a[10]), .B(n1873), .Z(n1420) );
  CENX1 U1948 ( .A(n1891), .B(n1408), .Z(n1135) );
  CND2X1 U1949 ( .A(n1421), .B(n1836), .Z(n44) );
  CND2X1 U1950 ( .A(n1416), .B(n82), .Z(n84) );
  CEOX1 U1951 ( .A(a[18]), .B(n1888), .Z(n1416) );
  CIVX1 U1952 ( .A(a[0]), .Z(n6) );
  CEOXL U1953 ( .A(a[20]), .B(n1891), .Z(n1415) );
  CND2X1 U1954 ( .A(n95), .B(n1414), .Z(n97) );
  CEOXL U1955 ( .A(a[22]), .B(n1894), .Z(n1414) );
  CNIVX1 U1956 ( .A(n116), .Z(n1898) );
  CND2X1 U1957 ( .A(n1622), .B(n333), .Z(n148) );
  CNIVX1 U1958 ( .A(n1402), .Z(n1841) );
  CNIVX1 U1959 ( .A(n1406), .Z(n1837) );
  CNIVX1 U1960 ( .A(n1404), .Z(n1839) );
  CNIVX1 U1961 ( .A(n116), .Z(n1899) );
  CNIVX1 U1962 ( .A(n1403), .Z(n1840) );
  CNIVX1 U1963 ( .A(n1401), .Z(n1842) );
  CND2X1 U1964 ( .A(n1825), .B(n1826), .Z(n1101) );
  CND2X1 U1965 ( .A(n1437), .B(n1824), .Z(n1826) );
  CND2X1 U1966 ( .A(n792), .B(n1642), .Z(n317) );
  COR2X1 U1967 ( .A(n792), .B(n1642), .Z(n1628) );
  CND2X1 U1968 ( .A(n1411), .B(n110), .Z(n112) );
  CEOXL U1969 ( .A(a[28]), .B(n109), .Z(n1411) );
  CEOX1 U1970 ( .A(n1852), .B(a[4]), .Z(n1629) );
  CIVX4 U1971 ( .A(n1629), .Z(n24) );
  CNIVX1 U1972 ( .A(n1405), .Z(n1838) );
  CND2X1 U1973 ( .A(n1410), .B(n114), .Z(n115) );
  CEOXL U1974 ( .A(n1816), .B(n147), .Z(n1901) );
  CND2XL U1975 ( .A(n365), .B(n1817), .Z(n147) );
  CENX1 U1976 ( .A(n1896), .B(n1839), .Z(n1107) );
  CENX1 U1977 ( .A(n1864), .B(n1838), .Z(n1279) );
  CENX1 U1978 ( .A(n1890), .B(n1838), .Z(n1132) );
  CENX1 U1979 ( .A(n1878), .B(n1838), .Z(n1183) );
  CENX1 U1980 ( .A(n1872), .B(n1838), .Z(n1227) );
  CENX1 U1981 ( .A(n1875), .B(n1838), .Z(n1204) );
  CENX1 U1982 ( .A(n1882), .B(n1838), .Z(n1164) );
  CND2XL U1983 ( .A(n1621), .B(n203), .Z(n126) );
  CNR2X1 U1984 ( .A(n214), .B(n1600), .Z(n196) );
  CENX1 U1985 ( .A(n1851), .B(n1389), .Z(n1323) );
  CENX1 U1986 ( .A(n1894), .B(n1407), .Z(n1121) );
  CND2X1 U1987 ( .A(n343), .B(n193), .Z(n125) );
  CIVX1 U1988 ( .A(n193), .Z(n191) );
  CENX1 U1989 ( .A(n1875), .B(n1844), .Z(n1198) );
  CENX1 U1990 ( .A(n1875), .B(n1843), .Z(n1199) );
  CIVX2 U1991 ( .A(n1407), .Z(n1824) );
  CENX1 U1992 ( .A(n1898), .B(n1887), .Z(n1151) );
  COND2XL U1993 ( .A(n69), .B(n1881), .C(n1188), .D(n66), .Z(n811) );
  CND2IX1 U1994 ( .B(n1899), .A(n1890), .Z(n1137) );
  CENX1 U1995 ( .A(n1883), .B(n1408), .Z(n1167) );
  CEO3X2 U1996 ( .A(n570), .B(n587), .C(n568), .Z(n564) );
  CND2X1 U1997 ( .A(n570), .B(n587), .Z(n1827) );
  CND2X1 U1998 ( .A(n570), .B(n568), .Z(n1828) );
  CND2XL U1999 ( .A(n587), .B(n568), .Z(n1829) );
  CND2XL U2000 ( .A(n566), .B(n585), .Z(n1830) );
  CND2X1 U2001 ( .A(n566), .B(n564), .Z(n1831) );
  CENX1 U2002 ( .A(n1891), .B(n1407), .Z(n1134) );
  COND2X1 U2003 ( .A(n91), .B(n1134), .C(n1133), .D(n89), .Z(n857) );
  CENX1 U2004 ( .A(n1862), .B(n1840), .Z(n1277) );
  CENX1 U2005 ( .A(n1862), .B(n1837), .Z(n1280) );
  CENX1 U2006 ( .A(n1896), .B(n1407), .Z(n1110) );
  CENX1 U2007 ( .A(n1875), .B(n1407), .Z(n1206) );
  CENX1 U2008 ( .A(n1883), .B(n1407), .Z(n1166) );
  CENX1 U2009 ( .A(n1879), .B(n1407), .Z(n1185) );
  CIVXL U2010 ( .A(n71), .Z(n1885) );
  CIVXL U2011 ( .A(n55), .Z(n1877) );
  CIVXL U2012 ( .A(n63), .Z(n1881) );
  CIVXL U2013 ( .A(n93), .Z(n1895) );
  CIVXL U2014 ( .A(n48), .Z(n1874) );
  CENX1 U2015 ( .A(n1896), .B(n1408), .Z(n1111) );
  CENX1 U2016 ( .A(n1879), .B(n1408), .Z(n1186) );
  CND2XL U2017 ( .A(n442), .B(n467), .Z(n1833) );
  CND2X1 U2018 ( .A(n442), .B(n444), .Z(n1834) );
  CND2XL U2019 ( .A(n467), .B(n444), .Z(n1835) );
  CND3XL U2020 ( .A(n1833), .B(n1834), .C(n1835), .Z(n439) );
  COND2X1 U2021 ( .A(n107), .B(n1437), .C(n105), .D(n1104), .Z(n805) );
  CEOXL U2022 ( .A(a[4]), .B(n1859), .Z(n1423) );
  CIVX1 U2023 ( .A(n226), .Z(n228) );
  CENX1 U2024 ( .A(n1861), .B(b[24]), .Z(n1259) );
  CENX1 U2025 ( .A(n1863), .B(a[8]), .Z(n42) );
  CND2XL U2026 ( .A(n340), .B(n172), .Z(n122) );
  CND2X1 U2027 ( .A(n440), .B(n465), .Z(n172) );
  CEOXL U2028 ( .A(n313), .B(n143), .Z(product[7]) );
  CEOXL U2029 ( .A(n321), .B(n145), .Z(n1900) );
  CNR2X1 U2030 ( .A(n171), .B(n176), .Z(n169) );
  CENX1 U2031 ( .A(n1856), .B(n1393), .Z(n1296) );
  CENXL U2032 ( .A(n1867), .B(n1393), .Z(n1240) );
  CENX1 U2033 ( .A(n1873), .B(n1393), .Z(n1215) );
  CENX1 U2034 ( .A(n1853), .B(n1392), .Z(n1326) );
  CENX1 U2035 ( .A(n1870), .B(n1392), .Z(n1239) );
  CENX1 U2036 ( .A(n1858), .B(n1392), .Z(n1295) );
  CEOXL U2037 ( .A(a[26]), .B(n104), .Z(n1412) );
  CIVXL U2038 ( .A(n21), .Z(n1860) );
  CND2X4 U2039 ( .A(n1420), .B(n50), .Z(n53) );
  CIVXL U2040 ( .A(n1854), .Z(n1850) );
  CIVXL U2041 ( .A(n1854), .Z(n1852) );
  CIVXL U2042 ( .A(n1854), .Z(n1853) );
  CIVXL U2043 ( .A(n1860), .Z(n1855) );
  CIVXL U2044 ( .A(n1860), .Z(n1856) );
  CIVXL U2045 ( .A(n1860), .Z(n1857) );
  CIVXL U2046 ( .A(n1860), .Z(n1858) );
  CIVXL U2047 ( .A(n1860), .Z(n1859) );
  CIVXL U2048 ( .A(n1866), .Z(n1862) );
  CIVXL U2049 ( .A(n1865), .Z(n1864) );
  CIVXL U2050 ( .A(n30), .Z(n1865) );
  CIVXL U2051 ( .A(n30), .Z(n1866) );
  CIVXL U2052 ( .A(n1871), .Z(n1867) );
  CIVXL U2053 ( .A(n1871), .Z(n1868) );
  CIVXL U2054 ( .A(n1871), .Z(n1869) );
  CIVXL U2055 ( .A(n1871), .Z(n1870) );
  CIVXL U2056 ( .A(n1881), .Z(n1878) );
  CIVXL U2057 ( .A(n1881), .Z(n1879) );
  CIVXL U2058 ( .A(n1881), .Z(n1880) );
  CIVXL U2059 ( .A(n1885), .Z(n1882) );
  CIVXL U2060 ( .A(n1885), .Z(n1883) );
  CIVXL U2061 ( .A(n1885), .Z(n1884) );
  CIVXL U2062 ( .A(n1889), .Z(n1886) );
  CIVXL U2063 ( .A(n1889), .Z(n1887) );
  CIVXL U2064 ( .A(n1889), .Z(n1888) );
  CIVXL U2065 ( .A(n79), .Z(n1889) );
  CIVXL U2066 ( .A(n1893), .Z(n1890) );
  CIVXL U2067 ( .A(n1893), .Z(n1891) );
  CIVXL U2068 ( .A(n1893), .Z(n1892) );
  CIVXL U2069 ( .A(n86), .Z(n1893) );
  CIVX2 U2070 ( .A(n1818), .Z(n365) );
  CIVX2 U2071 ( .A(n289), .Z(n357) );
  CIVX2 U2072 ( .A(n1582), .Z(n356) );
  CIVX2 U2073 ( .A(n275), .Z(n354) );
  CIVX2 U2074 ( .A(n248), .Z(n350) );
  CIVX2 U2075 ( .A(n171), .Z(n340) );
  CIVX2 U2076 ( .A(n333), .Z(n331) );
  CIVX2 U2077 ( .A(n1819), .Z(n323) );
  CIVX2 U2078 ( .A(n317), .Z(n315) );
  CIVX2 U2079 ( .A(n309), .Z(n307) );
  CIVX2 U2080 ( .A(n305), .Z(n304) );
  CIVX2 U2081 ( .A(n303), .Z(n301) );
  CIVX2 U2082 ( .A(n298), .Z(n296) );
  CIVX2 U2083 ( .A(n292), .Z(n291) );
  CIVX2 U2084 ( .A(n283), .Z(n282) );
  CIVX2 U2085 ( .A(n281), .Z(n279) );
  CIVX2 U2086 ( .A(n280), .Z(n355) );
  CIVX2 U2087 ( .A(n271), .Z(n269) );
  CIVX2 U2088 ( .A(n259), .Z(n261) );
  CIVX2 U2089 ( .A(n258), .Z(n352) );
  CIVX2 U2090 ( .A(n243), .Z(n241) );
  CIVX2 U2091 ( .A(n238), .Z(n236) );
  CIVX2 U2092 ( .A(n225), .Z(n347) );
  CIVX2 U2093 ( .A(n214), .Z(n216) );
  CIVX2 U2094 ( .A(n212), .Z(n210) );
  CIVX2 U2095 ( .A(n203), .Z(n201) );
  CIVX2 U2096 ( .A(n192), .Z(n343) );
  CIVX2 U2097 ( .A(n165), .Z(n163) );
  CIVX2 U2098 ( .A(n160), .Z(n158) );
  CIVX2 U2099 ( .A(n109), .Z(n1436) );
endmodule


module calc_DW02_mult_2_stage_4 ( A, B, TC, CLK, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC, CLK;
  wire   n15, n16, n17, \A_extended[32] , \B_extended[32] , n6, n8, n10, n11,
         n12, n13;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33;
  assign \A_extended[32]  = A[31];
  assign \B_extended[32]  = B[31];

  calc_DW_mult_tc_14 mult_96 ( .a({\A_extended[32] , \A_extended[32] , A[30:2], 
        1'b0, A[0]}), .b({\B_extended[32] , \B_extended[32] , B[30:0]}), 
        .product({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, PRODUCT[31:3], n15, 
        n16, n17}), .i_retiming_group_1_clk(CLK) );
  CFD1QXL clk_r_REG117_S1 ( .D(n16), .CP(CLK), .Q(n12) );
  CFD1QXL clk_r_REG194_S1 ( .D(n17), .CP(CLK), .Q(n11) );
  CFD1QXL clk_r_REG119_S1 ( .D(n15), .CP(CLK), .Q(n13) );
  CIVDXL U1 ( .A(n12), .Z1(n6) );
  CNIVX1 U2 ( .A(n6), .Z(PRODUCT[1]) );
  CIVDXL U3 ( .A(n11), .Z1(n8) );
  CNIVX1 U4 ( .A(n8), .Z(PRODUCT[0]) );
  CIVDXL U5 ( .A(n13), .Z1(n10) );
  CNIVX1 U6 ( .A(n10), .Z(PRODUCT[2]) );
endmodule


module calc_DW_mult_tc_15 ( a, b, product, i_retiming_group_1_clk );
  input [32:0] a;
  input [32:0] b;
  output [65:0] product;
  input i_retiming_group_1_clk;
  wire   n3, n9, n12, n15, n18, n21, n24, n27, n30, n33, n36, n39, n44, n48,
         n53, n55, n58, n61, n63, n66, n69, n71, n74, n77, n79, n82, n84, n86,
         n89, n91, n93, n95, n97, n99, n100, n102, n104, n105, n107, n109,
         n110, n112, n113, n114, n115, n116, n119, n121, n122, n123, n125,
         n126, n127, n128, n131, n132, n133, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n152, n154, n156, n158, n160, n163, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n179, n180, n181, n182,
         n184, n187, n188, n189, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n202, n203, n204, n205, n206, n210, n212, n213, n214,
         n215, n216, n217, n221, n223, n224, n225, n226, n228, n232, n233,
         n234, n236, n238, n239, n241, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n254, n256, n257, n258, n259, n261, n264,
         n265, n266, n267, n269, n271, n272, n273, n274, n275, n276, n277,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n296, n298, n299, n301, n303, n304,
         n305, n307, n309, n310, n311, n312, n313, n315, n317, n318, n319,
         n320, n321, n323, n325, n326, n327, n328, n329, n331, n333, n334,
         n335, n336, n340, n342, n343, n344, n347, n350, n352, n354, n355,
         n356, n357, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1410, n1411, n1412,
         n1413, n1414, n1415, n1417, n1419, n1422, n1424, n1435, n1436, n1437,
         n1438, n1439, n1440, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768;
  assign n3 = a[1];
  assign n12 = a[3];
  assign n21 = a[5];
  assign n30 = a[7];
  assign n39 = a[9];
  assign n48 = a[11];
  assign n55 = a[13];
  assign n63 = a[15];
  assign n71 = a[17];
  assign n79 = a[19];
  assign n86 = a[21];
  assign n93 = a[23];
  assign n99 = a[25];
  assign n104 = a[27];
  assign n109 = a[29];
  assign n113 = a[32];
  assign n116 = b[0];
  assign n1386 = b[23];
  assign n1387 = b[22];
  assign n1388 = b[21];
  assign n1389 = b[20];
  assign n1390 = b[19];
  assign n1391 = b[18];
  assign n1392 = b[17];
  assign n1393 = b[16];
  assign n1394 = b[15];
  assign n1395 = b[14];
  assign n1396 = b[13];
  assign n1397 = b[12];
  assign n1398 = b[11];
  assign n1399 = b[10];
  assign n1400 = b[9];
  assign n1401 = b[8];
  assign n1402 = b[7];
  assign n1403 = b[6];
  assign n1404 = b[5];
  assign n1405 = b[4];
  assign n1406 = b[3];
  assign n1407 = b[2];
  assign n1408 = b[1];
  assign n1685 = i_retiming_group_1_clk;

  CEO3X2 U375 ( .A(n387), .B(n369), .C(n385), .Z(n368) );
  CEO3X2 U376 ( .A(n1675), .B(n1677), .C(n1678), .Z(n369) );
  CEO3X2 U377 ( .A(n373), .B(n391), .C(n372), .Z(n370) );
  CEO3X2 U378 ( .A(n375), .B(n393), .C(n374), .Z(n371) );
  CEO3X2 U379 ( .A(n397), .B(n376), .C(n395), .Z(n372) );
  CEO3X2 U380 ( .A(n378), .B(n377), .C(n399), .Z(n373) );
  CEO3X2 U381 ( .A(n381), .B(n380), .C(n379), .Z(n374) );
  CEO3X2 U382 ( .A(n405), .B(n403), .C(n401), .Z(n375) );
  CEO3X2 U383 ( .A(n409), .B(n382), .C(n407), .Z(n376) );
  CEO3X2 U384 ( .A(n975), .B(n819), .C(n1029), .Z(n377) );
  CEO3X2 U385 ( .A(n891), .B(n951), .C(n1059), .Z(n378) );
  CEO3X2 U386 ( .A(n875), .B(n909), .C(n1001), .Z(n379) );
  CEO3X2 U387 ( .A(n803), .B(n849), .C(n929), .Z(n380) );
  CEO3X2 U388 ( .A(n831), .B(n821), .C(n861), .Z(n381) );
  CFA1X1 U390 ( .A(n388), .B(n386), .CI(n413), .CO(n383), .S(n384) );
  CFA1X1 U391 ( .A(n1673), .B(n1671), .CI(n1674), .CO(n385), .S(n386) );
  CFA1X1 U392 ( .A(n1672), .B(n1669), .CI(n1667), .CO(n387), .S(n388) );
  CFA1X1 U393 ( .A(n398), .B(n396), .CI(n421), .CO(n389), .S(n390) );
  CFA1X1 U394 ( .A(n425), .B(n400), .CI(n423), .CO(n391), .S(n392) );
  CFA1X1 U395 ( .A(n404), .B(n402), .CI(n427), .CO(n393), .S(n394) );
  CFA1X1 U396 ( .A(n410), .B(n406), .CI(n408), .CO(n395), .S(n396) );
  CFA1X1 U397 ( .A(n433), .B(n429), .CI(n431), .CO(n397), .S(n398) );
  CFA1X1 U398 ( .A(n1002), .B(n435), .CI(n437), .CO(n399), .S(n400) );
  CFA1X1 U399 ( .A(n910), .B(n1030), .CI(n976), .CO(n401), .S(n402) );
  CFA1X1 U400 ( .A(n892), .B(n1060), .CI(n930), .CO(n403), .S(n404) );
  CFA1X1 U402 ( .A(n822), .B(n862), .CI(n840), .CO(n407), .S(n408) );
  CFA1X1 U404 ( .A(n1670), .B(n414), .CI(n441), .CO(n411), .S(n412) );
  CFA1X1 U405 ( .A(n1666), .B(n1665), .CI(n1668), .CO(n413), .S(n414) );
  CFA1X1 U406 ( .A(n422), .B(n445), .CI(n447), .CO(n415), .S(n416) );
  CFA1X1 U407 ( .A(n426), .B(n424), .CI(n449), .CO(n417), .S(n418) );
  CFA1X1 U408 ( .A(n428), .B(n451), .CI(n453), .CO(n419), .S(n420) );
  CFA1X1 U409 ( .A(n434), .B(n430), .CI(n432), .CO(n421), .S(n422) );
  CFA1X1 U410 ( .A(n457), .B(n436), .CI(n455), .CO(n423), .S(n424) );
  CFA1X1 U411 ( .A(n463), .B(n459), .CI(n461), .CO(n425), .S(n426) );
  CFA1X1 U412 ( .A(n823), .B(n438), .CI(n1003), .CO(n427), .S(n428) );
  CFA1X1 U413 ( .A(n911), .B(n1031), .CI(n977), .CO(n429), .S(n430) );
  CFA1X1 U414 ( .A(n893), .B(n1061), .CI(n931), .CO(n431), .S(n432) );
  CFA1X1 U415 ( .A(n851), .B(n953), .CI(n877), .CO(n433), .S(n434) );
  CFA1X1 U416 ( .A(n833), .B(n863), .CI(n804), .CO(n435), .S(n436) );
  CHA1X1 U417 ( .A(n827), .B(n841), .CO(n437), .S(n438) );
  CFA1X1 U418 ( .A(n1664), .B(n442), .CI(n467), .CO(n439), .S(n440) );
  CFA1X1 U419 ( .A(n1662), .B(n1661), .CI(n1663), .CO(n441), .S(n442) );
  CFA1X1 U420 ( .A(n450), .B(n471), .CI(n473), .CO(n443), .S(n444) );
  CFA1X1 U421 ( .A(n454), .B(n452), .CI(n475), .CO(n445), .S(n446) );
  CFA1X1 U422 ( .A(n456), .B(n477), .CI(n479), .CO(n447), .S(n448) );
  CFA1X1 U423 ( .A(n462), .B(n458), .CI(n460), .CO(n449), .S(n450) );
  CFA1X1 U424 ( .A(n483), .B(n464), .CI(n481), .CO(n451), .S(n452) );
  CFA1X1 U425 ( .A(n489), .B(n485), .CI(n487), .CO(n453), .S(n454) );
  CFA1X1 U426 ( .A(n932), .B(n1032), .CI(n1004), .CO(n455), .S(n456) );
  CFA1X1 U427 ( .A(n912), .B(n1062), .CI(n954), .CO(n457), .S(n458) );
  CFA1X1 U428 ( .A(n864), .B(n978), .CI(n878), .CO(n459), .S(n460) );
  CFA1X1 U429 ( .A(n842), .B(n894), .CI(n852), .CO(n461), .S(n462) );
  CFA1X1 U430 ( .A(n824), .B(n1553), .CI(n828), .CO(n463), .S(n464) );
  CFA1X1 U431 ( .A(n1660), .B(n468), .CI(n1657), .CO(n465), .S(n466) );
  CFA1X1 U432 ( .A(n1658), .B(n1655), .CI(n1659), .CO(n467), .S(n468) );
  CFA1X1 U433 ( .A(n499), .B(n497), .CI(n476), .CO(n469), .S(n470) );
  CFA1X1 U434 ( .A(n480), .B(n478), .CI(n501), .CO(n471), .S(n472) );
  CFA1X1 U435 ( .A(n488), .B(n503), .CI(n482), .CO(n473), .S(n474) );
  CFA1X1 U437 ( .A(n507), .B(n511), .CI(n509), .CO(n477), .S(n478) );
  CFA1X1 U438 ( .A(n829), .B(n513), .CI(n490), .CO(n479), .S(n480) );
  CFA1X1 U439 ( .A(n1033), .B(n979), .CI(n1005), .CO(n481), .S(n482) );
  CFA1X1 U442 ( .A(n805), .B(n933), .CI(n865), .CO(n487), .S(n488) );
  CHA1X1 U443 ( .A(n835), .B(n843), .CO(n489), .S(n490) );
  CFA1X1 U444 ( .A(n1654), .B(n1656), .CI(n517), .CO(n491), .S(n492) );
  CFA1X1 U445 ( .A(n521), .B(n519), .CI(n498), .CO(n493), .S(n494) );
  CFA1X1 U446 ( .A(n523), .B(n500), .CI(n502), .CO(n495), .S(n496) );
  CFA1X1 U448 ( .A(n510), .B(n506), .CI(n508), .CO(n499), .S(n500) );
  CFA1X1 U449 ( .A(n529), .B(n512), .CI(n514), .CO(n501), .S(n502) );
  CFA1X1 U450 ( .A(n535), .B(n531), .CI(n533), .CO(n503), .S(n504) );
  CFA1X1 U453 ( .A(n866), .B(n980), .CI(n896), .CO(n509), .S(n510) );
  CFA1X1 U455 ( .A(n830), .B(n844), .CI(n836), .CO(n513), .S(n514) );
  CFA1X1 U456 ( .A(n1653), .B(n518), .CI(n1651), .CO(n515), .S(n516) );
  CFA1X1 U457 ( .A(n1647), .B(n1649), .CI(n1652), .CO(n517), .S(n518) );
  CFA1X1 U458 ( .A(n547), .B(n524), .CI(n526), .CO(n519), .S(n520) );
  CFA1X1 U459 ( .A(n551), .B(n528), .CI(n549), .CO(n521), .S(n522) );
  CFA1X1 U460 ( .A(n534), .B(n530), .CI(n532), .CO(n523), .S(n524) );
  CFA1X1 U461 ( .A(n555), .B(n536), .CI(n553), .CO(n525), .S(n526) );
  CFA1X1 U462 ( .A(n538), .B(n557), .CI(n559), .CO(n527), .S(n528) );
  CFA1X1 U463 ( .A(n981), .B(n1035), .CI(n837), .CO(n529), .S(n530) );
  CFA1X1 U464 ( .A(n957), .B(n1065), .CI(n897), .CO(n531), .S(n532) );
  CFA1X1 U466 ( .A(n935), .B(n806), .CI(n867), .CO(n535), .S(n536) );
  CHA1X1 U467 ( .A(n845), .B(n855), .CO(n537), .S(n538) );
  CFA1X1 U468 ( .A(n1648), .B(n1650), .CI(n1646), .CO(n539), .S(n540) );
  CFA1X1 U469 ( .A(n567), .B(n565), .CI(n546), .CO(n541), .S(n542) );
  CFA1X1 U470 ( .A(n569), .B(n548), .CI(n550), .CO(n543), .S(n544) );
  CFA1X1 U471 ( .A(n573), .B(n552), .CI(n571), .CO(n545), .S(n546) );
  CFA1X1 U472 ( .A(n556), .B(n554), .CI(n558), .CO(n547), .S(n548) );
  CFA1X1 U473 ( .A(n577), .B(n560), .CI(n575), .CO(n549), .S(n550) );
  CFA1X1 U474 ( .A(n1036), .B(n579), .CI(n581), .CO(n551), .S(n552) );
  CFA1X1 U475 ( .A(n916), .B(n1066), .CI(n958), .CO(n553), .S(n554) );
  CFA1X1 U476 ( .A(n882), .B(n936), .CI(n1574), .CO(n555), .S(n556) );
  CFA1X1 U478 ( .A(n838), .B(n856), .CI(n846), .CO(n559), .S(n560) );
  CFA1X1 U479 ( .A(n1644), .B(n1645), .CI(n1643), .CO(n561), .S(n562) );
  CFA1X1 U480 ( .A(n570), .B(n587), .CI(n568), .CO(n563), .S(n564) );
  CFA1X1 U481 ( .A(n591), .B(n589), .CI(n572), .CO(n565), .S(n566) );
  CFA1X1 U482 ( .A(n576), .B(n593), .CI(n574), .CO(n567), .S(n568) );
  CFA1X1 U483 ( .A(n595), .B(n578), .CI(n580), .CO(n569), .S(n570) );
  CFA1X1 U484 ( .A(n601), .B(n597), .CI(n599), .CO(n571), .S(n572) );
  CFA1X1 U485 ( .A(n1009), .B(n582), .CI(n1037), .CO(n573), .S(n574) );
  CFA1X1 U486 ( .A(n1548), .B(n983), .CI(n1067), .CO(n575), .S(n576) );
  CFA1X1 U487 ( .A(n869), .B(n847), .CI(n917), .CO(n577), .S(n578) );
  CFA1X1 U491 ( .A(n592), .B(n607), .CI(n590), .CO(n585), .S(n586) );
  CFA1X1 U492 ( .A(n611), .B(n609), .CI(n594), .CO(n587), .S(n588) );
  CFA1X1 U493 ( .A(n598), .B(n613), .CI(n596), .CO(n589), .S(n590) );
  CFA1X1 U494 ( .A(n615), .B(n600), .CI(n602), .CO(n591), .S(n592) );
  CFA1X1 U495 ( .A(n621), .B(n619), .CI(n617), .CO(n593), .S(n594) );
  CFA1X1 U496 ( .A(n918), .B(n1038), .CI(n984), .CO(n595), .S(n596) );
  CFA1X1 U497 ( .A(n900), .B(n1068), .CI(n960), .CO(n597), .S(n598) );
  CFA1X1 U498 ( .A(n884), .B(n1010), .CI(n938), .CO(n599), .S(n600) );
  CFA1X1 U499 ( .A(n848), .B(n858), .CI(n870), .CO(n601), .S(n602) );
  CFA1X1 U501 ( .A(n612), .B(n627), .CI(n610), .CO(n605), .S(n606) );
  CFA1X1 U502 ( .A(n631), .B(n629), .CI(n614), .CO(n607), .S(n608) );
  CFA1X1 U503 ( .A(n618), .B(n616), .CI(n633), .CO(n609), .S(n610) );
  CFA1X1 U504 ( .A(n635), .B(n620), .CI(n637), .CO(n611), .S(n612) );
  CFA1X1 U505 ( .A(n1039), .B(n639), .CI(n622), .CO(n613), .S(n614) );
  CFA1X1 U506 ( .A(n961), .B(n1069), .CI(n985), .CO(n615), .S(n616) );
  CFA1X1 U507 ( .A(n808), .B(n859), .CI(n901), .CO(n617), .S(n618) );
  CFA1X1 U508 ( .A(n885), .B(n1011), .CI(n939), .CO(n619), .S(n620) );
  CHA1X1 U509 ( .A(n871), .B(n919), .CO(n621), .S(n622) );
  CFA1X1 U510 ( .A(n1635), .B(n1636), .CI(n1634), .CO(n623), .S(n624) );
  CFA1X1 U511 ( .A(n632), .B(n645), .CI(n630), .CO(n625), .S(n626) );
  CFA1X1 U512 ( .A(n634), .B(n647), .CI(n649), .CO(n627), .S(n628) );
  CFA1X1 U513 ( .A(n638), .B(n640), .CI(n636), .CO(n629), .S(n630) );
  CFA1X1 U514 ( .A(n653), .B(n651), .CI(n655), .CO(n631), .S(n632) );
  CFA1X1 U515 ( .A(n986), .B(n657), .CI(n1012), .CO(n633), .S(n634) );
  CFA1X1 U517 ( .A(n902), .B(n1561), .CI(n1070), .CO(n637), .S(n638) );
  CFA1X1 U518 ( .A(n860), .B(n886), .CI(n872), .CO(n639), .S(n640) );
  CFA1X1 U519 ( .A(n1632), .B(n1633), .CI(n1631), .CO(n641), .S(n642) );
  CFA1X1 U520 ( .A(n650), .B(n663), .CI(n648), .CO(n643), .S(n644) );
  CFA1X1 U521 ( .A(n652), .B(n665), .CI(n667), .CO(n645), .S(n646) );
  CFA1X1 U522 ( .A(n669), .B(n654), .CI(n656), .CO(n647), .S(n648) );
  CFA1X1 U523 ( .A(n658), .B(n671), .CI(n673), .CO(n649), .S(n650) );
  CFA1X1 U524 ( .A(n987), .B(n1041), .CI(n873), .CO(n651), .S(n652) );
  CFA1X1 U525 ( .A(n903), .B(n1071), .CI(n921), .CO(n653), .S(n654) );
  CFA1X1 U526 ( .A(n809), .B(n1013), .CI(n941), .CO(n655), .S(n656) );
  CHA1X1 U527 ( .A(n887), .B(n963), .CO(n657), .S(n658) );
  CFA1X1 U528 ( .A(n1629), .B(n1630), .CI(n1628), .CO(n659), .S(n660) );
  CFA1X1 U529 ( .A(n668), .B(n679), .CI(n666), .CO(n661), .S(n662) );
  CFA1X1 U530 ( .A(n670), .B(n681), .CI(n683), .CO(n663), .S(n664) );
  CFA1X1 U531 ( .A(n685), .B(n672), .CI(n674), .CO(n665), .S(n666) );
  CFA1X1 U532 ( .A(n1014), .B(n687), .CI(n689), .CO(n667), .S(n668) );
  CFA1X1 U533 ( .A(n942), .B(n1042), .CI(n988), .CO(n669), .S(n670) );
  CFA1X1 U535 ( .A(n874), .B(n904), .CI(n888), .CO(n673), .S(n674) );
  CFA1X1 U536 ( .A(n1626), .B(n1627), .CI(n1625), .CO(n675), .S(n676) );
  CFA1X1 U537 ( .A(n684), .B(n695), .CI(n682), .CO(n677), .S(n678) );
  CFA1X1 U538 ( .A(n688), .B(n697), .CI(n686), .CO(n679), .S(n680) );
  CFA1X1 U539 ( .A(n703), .B(n699), .CI(n701), .CO(n681), .S(n682) );
  CFA1X1 U540 ( .A(n889), .B(n690), .CI(n1015), .CO(n683), .S(n684) );
  CFA1X1 U541 ( .A(n923), .B(n1043), .CI(n989), .CO(n685), .S(n686) );
  CFA1X1 U542 ( .A(n905), .B(n1073), .CI(n943), .CO(n687), .S(n688) );
  CHA1X1 U543 ( .A(n810), .B(n965), .CO(n689), .S(n690) );
  CFA1X1 U544 ( .A(n1623), .B(n1624), .CI(n1622), .CO(n691), .S(n692) );
  CFA1X1 U545 ( .A(n711), .B(n709), .CI(n698), .CO(n693), .S(n694) );
  CFA1X1 U546 ( .A(n704), .B(n700), .CI(n702), .CO(n695), .S(n696) );
  CFA1X1 U547 ( .A(n717), .B(n713), .CI(n715), .CO(n697), .S(n698) );
  CFA1X1 U548 ( .A(n966), .B(n1044), .CI(n1016), .CO(n699), .S(n700) );
  CFA1X1 U549 ( .A(n944), .B(n1074), .CI(n990), .CO(n701), .S(n702) );
  CFA1X1 U550 ( .A(n890), .B(n924), .CI(n906), .CO(n703), .S(n704) );
  CFA1X1 U551 ( .A(n1620), .B(n1621), .CI(n1617), .CO(n705), .S(n706) );
  CFA1X1 U552 ( .A(n714), .B(n712), .CI(n723), .CO(n707), .S(n708) );
  CFA1X1 U553 ( .A(n727), .B(n725), .CI(n716), .CO(n709), .S(n710) );
  CFA1X1 U554 ( .A(n907), .B(n729), .CI(n718), .CO(n711), .S(n712) );
  CFA1X1 U555 ( .A(n991), .B(n1045), .CI(n1017), .CO(n713), .S(n714) );
  CFA1X1 U556 ( .A(n925), .B(n1075), .CI(n945), .CO(n715), .S(n716) );
  CHA1X1 U557 ( .A(n811), .B(n967), .CO(n717), .S(n718) );
  CFA1X1 U558 ( .A(n724), .B(n722), .CI(n733), .CO(n719), .S(n720) );
  CFA1X1 U559 ( .A(n728), .B(n735), .CI(n726), .CO(n721), .S(n722) );
  CFA1X1 U560 ( .A(n739), .B(n730), .CI(n737), .CO(n723), .S(n724) );
  CFA1X1 U564 ( .A(n736), .B(n734), .CI(n745), .CO(n731), .S(n732) );
  CFA1X1 U565 ( .A(n740), .B(n747), .CI(n738), .CO(n733), .S(n734) );
  CFA1X1 U566 ( .A(n742), .B(n749), .CI(n751), .CO(n735), .S(n736) );
  CFA1X1 U567 ( .A(n969), .B(n1047), .CI(n1019), .CO(n737), .S(n738) );
  CFA1X1 U570 ( .A(n755), .B(n746), .CI(n748), .CO(n743), .S(n744) );
  CFA1X1 U571 ( .A(n752), .B(n757), .CI(n750), .CO(n745), .S(n746) );
  CFA1X1 U572 ( .A(n1020), .B(n759), .CI(n761), .CO(n747), .S(n748) );
  CFA1X1 U573 ( .A(n1078), .B(n994), .CI(n1048), .CO(n749), .S(n750) );
  CFA1X1 U574 ( .A(n928), .B(n970), .CI(n948), .CO(n751), .S(n752) );
  CFA1X1 U575 ( .A(n758), .B(n756), .CI(n765), .CO(n753), .S(n754) );
  CFA1X1 U576 ( .A(n769), .B(n760), .CI(n767), .CO(n755), .S(n756) );
  CFA1X1 U577 ( .A(n995), .B(n762), .CI(n1049), .CO(n757), .S(n758) );
  CFA1X1 U578 ( .A(n971), .B(n1079), .CI(n1021), .CO(n759), .S(n760) );
  CHA1X1 U579 ( .A(n813), .B(n949), .CO(n761), .S(n762) );
  CFA1X1 U580 ( .A(n768), .B(n766), .CI(n773), .CO(n763), .S(n764) );
  CFA1X1 U581 ( .A(n777), .B(n770), .CI(n775), .CO(n765), .S(n766) );
  CFA1X1 U582 ( .A(n1022), .B(n1080), .CI(n1050), .CO(n767), .S(n768) );
  CFA1X1 U583 ( .A(n950), .B(n1565), .CI(n972), .CO(n769), .S(n770) );
  CFA1X1 U584 ( .A(n781), .B(n774), .CI(n776), .CO(n771), .S(n772) );
  CFA1X1 U585 ( .A(n973), .B(n783), .CI(n778), .CO(n773), .S(n774) );
  CFA1X1 U586 ( .A(n997), .B(n1081), .CI(n1023), .CO(n775), .S(n776) );
  CHA1X1 U587 ( .A(n814), .B(n1051), .CO(n777), .S(n778) );
  CFA1X1 U588 ( .A(n787), .B(n782), .CI(n784), .CO(n779), .S(n780) );
  CFA1X1 U589 ( .A(n1052), .B(n789), .CI(n1082), .CO(n781), .S(n782) );
  CFA1X1 U590 ( .A(n974), .B(n1024), .CI(n998), .CO(n783), .S(n784) );
  CFA1X1 U591 ( .A(n790), .B(n788), .CI(n793), .CO(n785), .S(n786) );
  CHA1X1 U593 ( .A(n815), .B(n999), .CO(n789), .S(n790) );
  CFA1X1 U594 ( .A(n1084), .B(n794), .CI(n797), .CO(n791), .S(n792) );
  CFA1X1 U596 ( .A(n1055), .B(n798), .CI(n1085), .CO(n795), .S(n796) );
  CHA1X1 U597 ( .A(n816), .B(n1027), .CO(n797), .S(n798) );
  CFA1X1 U598 ( .A(n1028), .B(n1086), .CI(n1056), .CO(n799), .S(n800) );
  CHA1X1 U599 ( .A(n817), .B(n1087), .CO(n801), .S(n802) );
  COND2X1 U600 ( .A(n1092), .B(n114), .C(n1435), .D(n115), .Z(n803) );
  COND2X1 U601 ( .A(n1091), .B(n115), .C(n114), .D(n1090), .Z(n819) );
  CND2IX1 U605 ( .B(n1710), .A(n113), .Z(n1092) );
  COND2X1 U606 ( .A(n1097), .B(n110), .C(n1436), .D(n112), .Z(n804) );
  COND2X1 U608 ( .A(n112), .B(n1095), .C(n110), .D(n1094), .Z(n822) );
  CND2IX1 U615 ( .B(n1710), .A(n109), .Z(n1097) );
  COND2X1 U620 ( .A(n107), .B(n1102), .C(n105), .D(n1101), .Z(n828) );
  CND2IX1 U629 ( .B(n1710), .A(n104), .Z(n1104) );
  COND2X1 U636 ( .A(n1552), .B(n1111), .C(n100), .D(n1110), .Z(n836) );
  COND2X1 U637 ( .A(n1112), .B(n1552), .C(n100), .D(n1111), .Z(n837) );
  CND2IX1 U647 ( .B(n1710), .A(n1708), .Z(n1113) );
  COND2X1 U670 ( .A(n91), .B(n1440), .C(n89), .D(n1137), .Z(n808) );
  COND2X1 U671 ( .A(n91), .B(n1126), .C(n1125), .D(n89), .Z(n849) );
  COND2X1 U672 ( .A(n91), .B(n1127), .C(n1126), .D(n89), .Z(n850) );
  COND2X1 U673 ( .A(n91), .B(n1128), .C(n1127), .D(n89), .Z(n851) );
  COND2X1 U674 ( .A(n91), .B(n1129), .C(n1128), .D(n89), .Z(n852) );
  COND2X1 U675 ( .A(n91), .B(n1130), .C(n1129), .D(n89), .Z(n853) );
  COND2X1 U676 ( .A(n91), .B(n1131), .C(n1130), .D(n89), .Z(n854) );
  COND2X1 U677 ( .A(n91), .B(n1132), .C(n1131), .D(n89), .Z(n855) );
  COND2X1 U678 ( .A(n91), .B(n1133), .C(n1132), .D(n89), .Z(n856) );
  COND2X1 U680 ( .A(n91), .B(n1135), .C(n1134), .D(n89), .Z(n858) );
  COND2X1 U681 ( .A(n1136), .B(n91), .C(n89), .D(n1135), .Z(n859) );
  COND2X1 U696 ( .A(n84), .B(n1767), .C(n82), .D(n1152), .Z(n809) );
  COND2X1 U699 ( .A(n84), .B(n1141), .C(n1140), .D(n82), .Z(n863) );
  COND2X1 U700 ( .A(n84), .B(n1142), .C(n1141), .D(n82), .Z(n864) );
  COND2X1 U702 ( .A(n84), .B(n1144), .C(n1143), .D(n82), .Z(n866) );
  COND2X1 U704 ( .A(n84), .B(n1146), .C(n1145), .D(n82), .Z(n868) );
  COND2X1 U706 ( .A(n84), .B(n1148), .C(n1147), .D(n82), .Z(n870) );
  COND2X1 U707 ( .A(n84), .B(n1149), .C(n1148), .D(n82), .Z(n871) );
  COND2X1 U708 ( .A(n84), .B(n1150), .C(n1149), .D(n82), .Z(n872) );
  CND2IX1 U725 ( .B(n1710), .A(n1763), .Z(n1152) );
  CND2IX1 U759 ( .B(n1710), .A(n1686), .Z(n1169) );
  COND2X1 U766 ( .A(n69), .B(n1176), .C(n1175), .D(n66), .Z(n896) );
  COND2X1 U767 ( .A(n69), .B(n1177), .C(n1176), .D(n66), .Z(n897) );
  COND2X1 U770 ( .A(n69), .B(n1180), .C(n1179), .D(n66), .Z(n900) );
  COND2X1 U771 ( .A(n69), .B(n1181), .C(n1180), .D(n66), .Z(n901) );
  COND2X1 U773 ( .A(n69), .B(n1183), .C(n1182), .D(n66), .Z(n903) );
  COND2X1 U774 ( .A(n69), .B(n1184), .C(n1183), .D(n66), .Z(n904) );
  COND2X1 U776 ( .A(n69), .B(n1186), .C(n1185), .D(n66), .Z(n906) );
  COND2X1 U803 ( .A(n61), .B(n1194), .C(n1193), .D(n1549), .Z(n913) );
  COND2X1 U805 ( .A(n61), .B(n1196), .C(n1195), .D(n1550), .Z(n915) );
  COND2X1 U806 ( .A(n61), .B(n1197), .C(n1196), .D(n1550), .Z(n916) );
  COND2X1 U809 ( .A(n61), .B(n1200), .C(n1199), .D(n1550), .Z(n919) );
  COND2X1 U847 ( .A(n53), .B(n1217), .C(n1216), .D(n1583), .Z(n935) );
  COND2X1 U851 ( .A(n53), .B(n1221), .C(n1220), .D(n1583), .Z(n939) );
  COND2X1 U893 ( .A(n44), .B(n1240), .C(n1239), .D(n1582), .Z(n957) );
  COND2X1 U894 ( .A(n44), .B(n1241), .C(n1240), .D(n1582), .Z(n958) );
  COND2X1 U895 ( .A(n44), .B(n1242), .C(n1241), .D(n1582), .Z(n959) );
  COND2X1 U896 ( .A(n44), .B(n1243), .C(n1242), .D(n1582), .Z(n960) );
  COND2X1 U897 ( .A(n44), .B(n1244), .C(n1243), .D(n1582), .Z(n961) );
  COND2X1 U908 ( .A(n44), .B(n1255), .C(n1254), .D(n1582), .Z(n972) );
  CND2IX1 U935 ( .B(n1710), .A(n1740), .Z(n1257) );
  COND2X1 U943 ( .A(n36), .B(n1265), .C(n1264), .D(n33), .Z(n981) );
  COND2X1 U944 ( .A(n36), .B(n1266), .C(n1265), .D(n33), .Z(n982) );
  COND2X1 U1051 ( .A(n18), .B(n1317), .C(n1316), .D(n15), .Z(n1031) );
  COND2X1 U1053 ( .A(n18), .B(n1319), .C(n1318), .D(n15), .Z(n1033) );
  COND2X1 U1056 ( .A(n18), .B(n1322), .C(n1321), .D(n15), .Z(n1036) );
  COND2X1 U1057 ( .A(n18), .B(n1323), .C(n1322), .D(n15), .Z(n1037) );
  COND2X1 U1058 ( .A(n18), .B(n1324), .C(n1323), .D(n15), .Z(n1038) );
  COND2X1 U1060 ( .A(n18), .B(n1326), .C(n1325), .D(n15), .Z(n1040) );
  COND2X1 U1062 ( .A(n18), .B(n1328), .C(n1327), .D(n15), .Z(n1042) );
  COND2X1 U1063 ( .A(n18), .B(n1329), .C(n1328), .D(n15), .Z(n1043) );
  COND2X1 U1064 ( .A(n18), .B(n1330), .C(n1329), .D(n15), .Z(n1044) );
  COND2X1 U1065 ( .A(n18), .B(n1331), .C(n1330), .D(n15), .Z(n1045) );
  COND2X1 U1067 ( .A(n18), .B(n1333), .C(n1332), .D(n15), .Z(n1047) );
  COND2X1 U1068 ( .A(n18), .B(n1334), .C(n1333), .D(n15), .Z(n1048) );
  COND2X1 U1076 ( .A(n18), .B(n1342), .C(n1341), .D(n15), .Z(n1056) );
  COND2X1 U1110 ( .A(n9), .B(n1718), .C(n1713), .D(n1377), .Z(n818) );
  COND2X1 U1111 ( .A(n9), .B(n1346), .C(n1713), .D(n1345), .Z(n1059) );
  COND2X1 U1112 ( .A(n9), .B(n1347), .C(n1713), .D(n1346), .Z(n1060) );
  COND2X1 U1113 ( .A(n9), .B(n1348), .C(n1713), .D(n1347), .Z(n1061) );
  COND2X1 U1114 ( .A(n9), .B(n1349), .C(n1713), .D(n1348), .Z(n1062) );
  COND2X1 U1115 ( .A(n9), .B(n1350), .C(n1713), .D(n1349), .Z(n1063) );
  COND2X1 U1116 ( .A(n9), .B(n1351), .C(n1713), .D(n1350), .Z(n1064) );
  COND2X1 U1117 ( .A(n9), .B(n1352), .C(n1713), .D(n1351), .Z(n1065) );
  COND2X1 U1118 ( .A(n9), .B(n1353), .C(n1713), .D(n1352), .Z(n1066) );
  COND2X1 U1119 ( .A(n9), .B(n1354), .C(n1713), .D(n1353), .Z(n1067) );
  COND2X1 U1120 ( .A(n9), .B(n1355), .C(n1713), .D(n1354), .Z(n1068) );
  COND2X1 U1121 ( .A(n9), .B(n1356), .C(n1713), .D(n1355), .Z(n1069) );
  COND2X1 U1122 ( .A(n9), .B(n1357), .C(n1714), .D(n1356), .Z(n1070) );
  COND2X1 U1123 ( .A(n9), .B(n1358), .C(n1714), .D(n1357), .Z(n1071) );
  COND2X1 U1124 ( .A(n9), .B(n1359), .C(n1714), .D(n1358), .Z(n1072) );
  COND2X1 U1125 ( .A(n9), .B(n1360), .C(n1714), .D(n1359), .Z(n1073) );
  COND2X1 U1126 ( .A(n9), .B(n1361), .C(n1713), .D(n1360), .Z(n1074) );
  COND2X1 U1127 ( .A(n9), .B(n1362), .C(n1713), .D(n1361), .Z(n1075) );
  COND2X1 U1128 ( .A(n9), .B(n1363), .C(n1713), .D(n1362), .Z(n1076) );
  COND2X1 U1129 ( .A(n9), .B(n1364), .C(n1713), .D(n1363), .Z(n1077) );
  COND2X1 U1130 ( .A(n9), .B(n1365), .C(n1713), .D(n1364), .Z(n1078) );
  COND2X1 U1131 ( .A(n9), .B(n1366), .C(n1713), .D(n1365), .Z(n1079) );
  COND2X1 U1132 ( .A(n9), .B(n1367), .C(n1713), .D(n1366), .Z(n1080) );
  COND2X1 U1133 ( .A(n9), .B(n1368), .C(n1713), .D(n1367), .Z(n1081) );
  COND2X1 U1134 ( .A(n9), .B(n1369), .C(n1713), .D(n1368), .Z(n1082) );
  COND2X1 U1135 ( .A(n9), .B(n1370), .C(n1713), .D(n1369), .Z(n1083) );
  COND2X1 U1136 ( .A(n9), .B(n1371), .C(n1713), .D(n1370), .Z(n1084) );
  COND2X1 U1137 ( .A(n9), .B(n1372), .C(n1713), .D(n1371), .Z(n1085) );
  COND2X1 U1138 ( .A(n9), .B(n1373), .C(n1713), .D(n1372), .Z(n1086) );
  COND2X1 U1139 ( .A(n9), .B(n1374), .C(n1713), .D(n1373), .Z(n1087) );
  COND2X1 U1140 ( .A(n9), .B(n1375), .C(n1713), .D(n1374), .Z(n1088) );
  COND2X1 U1141 ( .A(n9), .B(n1376), .C(n1713), .D(n1375), .Z(n1089) );
  CFD1QXL clk_r_REG232_S1 ( .D(n389), .CP(n1685), .Q(n1675) );
  CFD1QXL clk_r_REG217_S1 ( .D(n370), .CP(n1685), .Q(n1678) );
  CFD1QXL clk_r_REG198_S1 ( .D(n443), .CP(n1685), .Q(n1665) );
  CFD1QXL clk_r_REG201_S1 ( .D(n415), .CP(n1685), .Q(n1671) );
  CFD1QXL clk_r_REG215_S1 ( .D(n542), .CP(n1685), .Q(n1650) );
  CFD1QXL clk_r_REG206_S1 ( .D(n469), .CP(n1685), .Q(n1661) );
  CFD1QXL clk_r_REG205_S1 ( .D(n494), .CP(n1685), .Q(n1656) );
  CFD1QXL clk_r_REG210_S1 ( .D(n564), .CP(n1685), .Q(n1645) );
  CFD1QXL clk_r_REG224_S1 ( .D(n287), .CP(n1685), .Q(n1681) );
  CFD1QXL clk_r_REG264_S1 ( .D(n418), .CP(n1685), .Q(n1668) );
  CFD1QXL clk_r_REG233_S1 ( .D(n390), .CP(n1685), .Q(n1674) );
  CFD1QXL clk_r_REG261_S1 ( .D(n419), .CP(n1685), .Q(n1667) );
  CFD1QXL clk_r_REG209_S1 ( .D(n563), .CP(n1685), .Q(n1646) );
  CFD1QXL clk_r_REG204_S1 ( .D(n493), .CP(n1685), .Q(n1657) );
  CFD1QXL clk_r_REG214_S1 ( .D(n541), .CP(n1685), .Q(n1651) );
  CFD1QXL clk_r_REG256_S1 ( .D(n585), .CP(n1685), .Q(n1643) );
  CFD1QXL clk_r_REG262_S1 ( .D(n420), .CP(n1685), .Q(n1666) );
  CFD1QXL clk_r_REG269_S1 ( .D(n394), .CP(n1685), .Q(n1672) );
  CFD1QXL clk_r_REG199_S1 ( .D(n444), .CP(n1685), .Q(n1664) );
  CFD1QXL clk_r_REG202_S1 ( .D(n416), .CP(n1685), .Q(n1670) );
  CFD1QXL clk_r_REG212_S1 ( .D(n544), .CP(n1685), .Q(n1648) );
  CFD1QXL clk_r_REG207_S1 ( .D(n470), .CP(n1685), .Q(n1660) );
  CFD1QXL clk_r_REG196_S1 ( .D(n496), .CP(n1685), .Q(n1654) );
  CFD1QXL clk_r_REG267_S1 ( .D(n305), .CP(n1685), .Q(n1676) );
  CFD1QXL clk_r_REG228_S1 ( .D(n732), .CP(n1685), .Q(n1615) );
  CFD1QXL clk_r_REG238_S1 ( .D(n625), .CP(n1685), .Q(n1637) );
  CFD1QXL clk_r_REG243_S1 ( .D(n605), .CP(n1685), .Q(n1640) );
  CFD1QXL clk_r_REG225_S1 ( .D(n286), .CP(n1685), .Q(n1682) );
  CFD1QXL clk_r_REG257_S1 ( .D(n586), .CP(n1685), .Q(n1642) );
  CFD1QXL clk_r_REG244_S1 ( .D(n606), .CP(n1685), .Q(n1639) );
  CFD1QXL clk_r_REG219_S1 ( .D(n1595), .CP(n1685), .Q(n1683) );
  CFD1QXL clk_r_REG255_S1 ( .D(n608), .CP(n1685), .Q(n1638) );
  CFD1QXL clk_r_REG258_S1 ( .D(n588), .CP(n1685), .Q(n1641) );
  CFD1QXL clk_r_REG236_S1 ( .D(n662), .CP(n1685), .Q(n1630) );
  CFD1QXL clk_r_REG239_S1 ( .D(n626), .CP(n1685), .Q(n1636) );
  CFD1QXL clk_r_REG241_S1 ( .D(n644), .CP(n1685), .Q(n1633) );
  CFD1QXL clk_r_REG240_S1 ( .D(n643), .CP(n1685), .Q(n1634) );
  CFD1QXL clk_r_REG235_S1 ( .D(n661), .CP(n1685), .Q(n1631) );
  CFD1QXL clk_r_REG242_S1 ( .D(n628), .CP(n1685), .Q(n1635) );
  CFD1QXL clk_r_REG237_S1 ( .D(n646), .CP(n1685), .Q(n1632) );
  CFD1QXL clk_r_REG220_S1 ( .D(n298), .CP(n1685), .Q(n1680) );
  CFD1QXL clk_r_REG218_S1 ( .D(n303), .CP(n1685), .Q(n1679) );
  CFD1QXL clk_r_REG223_S1 ( .D(n754), .CP(n1685), .Q(n1613) );
  CFD1QXL clk_r_REG230_S1 ( .D(n719), .CP(n1685), .Q(n1619) );
  CFD1QXL clk_r_REG222_S1 ( .D(n763), .CP(n1685), .Q(n1612) );
  CFD1QXL clk_r_REG221_S1 ( .D(n1594), .CP(n1685), .Q(n1684) );
  CFD1QXL clk_r_REG231_S1 ( .D(n720), .CP(n1685), .Q(n1618) );
  CFD1QXL clk_r_REG227_S1 ( .D(n731), .CP(n1685), .Q(n1616) );
  CFD1QX2 clk_r_REG254_S1 ( .D(n710), .CP(n1685), .Q(n1620) );
  CFD1QX1 clk_r_REG229_S1 ( .D(n721), .CP(n1685), .Q(n1617) );
  CFD1QX1 clk_r_REG253_S1 ( .D(n696), .CP(n1685), .Q(n1623) );
  CFD1QX1 clk_r_REG252_S1 ( .D(n680), .CP(n1685), .Q(n1626) );
  CFD1QX1 clk_r_REG250_S1 ( .D(n693), .CP(n1685), .Q(n1625) );
  CFD1QX2 clk_r_REG200_S1 ( .D(n448), .CP(n1685), .Q(n1662) );
  CFD1QX1 clk_r_REG208_S1 ( .D(n474), .CP(n1685), .Q(n1658) );
  CFD1QX1 clk_r_REG248_S1 ( .D(n707), .CP(n1685), .Q(n1622) );
  CFD1QX2 clk_r_REG249_S1 ( .D(n708), .CP(n1685), .Q(n1621) );
  CFD1QX1 clk_r_REG213_S1 ( .D(n545), .CP(n1685), .Q(n1647) );
  CFD1QX2 clk_r_REG246_S1 ( .D(n678), .CP(n1685), .Q(n1627) );
  CFD1QX2 clk_r_REG216_S1 ( .D(n522), .CP(n1685), .Q(n1652) );
  CFD1QX1 clk_r_REG247_S1 ( .D(n664), .CP(n1685), .Q(n1629) );
  CFD1QX2 clk_r_REG197_S1 ( .D(n472), .CP(n1685), .Q(n1659) );
  CFD1QX2 clk_r_REG251_S1 ( .D(n694), .CP(n1685), .Q(n1624) );
  CFD1QX1 clk_r_REG260_S1 ( .D(n446), .CP(n1685), .Q(n1663) );
  CFD1QX1 clk_r_REG245_S1 ( .D(n677), .CP(n1685), .Q(n1628) );
  CFD1QX2 clk_r_REG259_S1 ( .D(n566), .CP(n1685), .Q(n1644) );
  CFD1QXL clk_r_REG234_S1 ( .D(n371), .CP(n1685), .Q(n1677) );
  CFD1QXL clk_r_REG265_S1 ( .D(n392), .CP(n1685), .Q(n1673) );
  CFD1QXL clk_r_REG203_S1 ( .D(n520), .CP(n1685), .Q(n1653) );
  CFD1QXL clk_r_REG263_S1 ( .D(n417), .CP(n1685), .Q(n1669) );
  CFD1QXL clk_r_REG226_S1 ( .D(n743), .CP(n1685), .Q(n1614) );
  CFD1QX1 clk_r_REG195_S1 ( .D(n495), .CP(n1685), .Q(n1655) );
  CFD1QX1 clk_r_REG211_S1 ( .D(n543), .CP(n1685), .Q(n1649) );
  COND1X1 U1271 ( .A(n205), .B(n1567), .C(n206), .Z(n204) );
  CENXL U1272 ( .A(n250), .B(n132), .Z(product[18]) );
  CFA1XL U1273 ( .A(n947), .B(n1077), .CI(n993), .CO(n739), .S(n740) );
  CIVX1 U1274 ( .A(n937), .Z(n1547) );
  CIVX2 U1275 ( .A(n1547), .Z(n1548) );
  COND2XL U1276 ( .A(n27), .B(n1306), .C(n1305), .D(n24), .Z(n1021) );
  CENX2 U1277 ( .A(a[14]), .B(n1754), .Z(n1588) );
  CENX2 U1278 ( .A(n1748), .B(a[12]), .Z(n1549) );
  CENX2 U1279 ( .A(n1748), .B(a[12]), .Z(n1550) );
  CENX2 U1280 ( .A(n1748), .B(a[12]), .Z(n58) );
  COND2X2 U1281 ( .A(n1104), .B(n105), .C(n1437), .D(n107), .Z(n805) );
  CENX2 U1282 ( .A(n1708), .B(a[26]), .Z(n105) );
  CENX1 U1283 ( .A(n1551), .B(n1708), .Z(n1413) );
  CIVX20 U1284 ( .A(a[24]), .Z(n1551) );
  CND2X2 U1285 ( .A(n1413), .B(n100), .Z(n1552) );
  CND2X1 U1286 ( .A(n1413), .B(n100), .Z(n102) );
  COND2XL U1287 ( .A(n84), .B(n1139), .C(n1138), .D(n82), .Z(n861) );
  CENXL U1288 ( .A(n1766), .B(n1396), .Z(n1138) );
  COND2XL U1289 ( .A(n84), .B(n1140), .C(n1139), .D(n82), .Z(n862) );
  COND2XL U1290 ( .A(n1151), .B(n84), .C(n82), .D(n1150), .Z(n873) );
  COND2XL U1291 ( .A(n84), .B(n1147), .C(n1146), .D(n82), .Z(n869) );
  CENXL U1292 ( .A(n1709), .B(n1766), .Z(n1151) );
  CENXL U1293 ( .A(n1711), .B(n1766), .Z(n1150) );
  COND2X1 U1294 ( .A(n107), .B(n1100), .C(n105), .D(n1099), .Z(n826) );
  COND2XL U1295 ( .A(n107), .B(n1099), .C(n105), .D(n1098), .Z(n825) );
  COND2XL U1296 ( .A(n107), .B(n1101), .C(n105), .D(n1100), .Z(n827) );
  COND2X1 U1297 ( .A(n1103), .B(n107), .C(n105), .D(n1102), .Z(n829) );
  COND2X1 U1298 ( .A(n18), .B(n1321), .C(n1320), .D(n15), .Z(n1035) );
  CENX2 U1299 ( .A(a[0]), .B(n1717), .Z(n1587) );
  CIVX4 U1300 ( .A(n1585), .Z(n9) );
  CFA1XL U1301 ( .A(n914), .B(n1064), .CI(n934), .CO(n507), .S(n508) );
  CFA1X1 U1302 ( .A(n895), .B(n1063), .CI(n913), .CO(n483), .S(n484) );
  COND2X1 U1303 ( .A(n69), .B(n1175), .C(n1174), .D(n66), .Z(n895) );
  CNIVX1 U1304 ( .A(n834), .Z(n1553) );
  COND1X2 U1305 ( .A(n193), .B(n187), .C(n188), .Z(n182) );
  CIVX2 U1306 ( .A(n21), .Z(n1733) );
  CND2XL U1307 ( .A(n1411), .B(n110), .Z(n112) );
  COND2X1 U1308 ( .A(n1113), .B(n100), .C(n1438), .D(n102), .Z(n806) );
  CNR2IXL U1309 ( .B(n1710), .A(n100), .Z(n838) );
  CND2IX2 U1310 ( .B(n1584), .A(n1582), .Z(n44) );
  CANR1X1 U1311 ( .A(n181), .B(n194), .C(n182), .Z(n180) );
  CIVX2 U1312 ( .A(n30), .Z(n1739) );
  CIVX2 U1313 ( .A(n1739), .Z(n1735) );
  CIVX1 U1314 ( .A(n39), .Z(n1746) );
  CIVX2 U1315 ( .A(a[0]), .Z(n1714) );
  CIVX2 U1316 ( .A(a[0]), .Z(n1713) );
  CIVX1 U1317 ( .A(n30), .Z(n1738) );
  CIVDXL U1318 ( .A(n176), .Z0(n1554), .Z1(n1555) );
  CAN2XL U1319 ( .A(n1605), .B(n1603), .Z(n1556) );
  COND2X1 U1320 ( .A(n91), .B(n1134), .C(n1133), .D(n89), .Z(n857) );
  CNR2X2 U1321 ( .A(n466), .B(n491), .Z(n176) );
  COND2XL U1322 ( .A(n44), .B(n1249), .C(n1248), .D(n1582), .Z(n966) );
  COND2XL U1323 ( .A(n44), .B(n1238), .C(n1237), .D(n1582), .Z(n955) );
  COND2XL U1324 ( .A(n44), .B(n1247), .C(n1246), .D(n1582), .Z(n964) );
  COND2XL U1325 ( .A(n44), .B(n1254), .C(n1253), .D(n1582), .Z(n971) );
  COND2XL U1326 ( .A(n44), .B(n1239), .C(n1238), .D(n1582), .Z(n956) );
  CENXL U1327 ( .A(n1722), .B(n1700), .Z(n1341) );
  CENXL U1328 ( .A(n1722), .B(n1706), .Z(n1338) );
  CENXL U1329 ( .A(n1722), .B(n1702), .Z(n1340) );
  CENXL U1330 ( .A(n1722), .B(n1704), .Z(n1339) );
  CENXL U1331 ( .A(n1709), .B(n1744), .Z(n1256) );
  CND2X4 U1332 ( .A(n1417), .B(n74), .Z(n77) );
  CEOX2 U1333 ( .A(a[16]), .B(n1590), .Z(n1417) );
  CEOX2 U1334 ( .A(a[22]), .B(n1707), .Z(n1414) );
  CNIVX4 U1335 ( .A(n93), .Z(n1707) );
  CENX1 U1336 ( .A(n504), .B(n1557), .Z(n498) );
  CENX1 U1337 ( .A(n527), .B(n525), .Z(n1557) );
  CIVXL U1338 ( .A(n920), .Z(n1558) );
  CIVX2 U1339 ( .A(n1558), .Z(n1559) );
  CFA1X1 U1340 ( .A(n1559), .B(n1040), .CI(n940), .CO(n635), .S(n636) );
  CND2X1 U1341 ( .A(n344), .B(n1602), .Z(n198) );
  CENX1 U1342 ( .A(n224), .B(n128), .Z(product[22]) );
  COND1X1 U1343 ( .A(n225), .B(n1567), .C(n226), .Z(n224) );
  COND2X1 U1344 ( .A(n53), .B(n1222), .C(n1221), .D(n1583), .Z(n940) );
  CENX4 U1345 ( .A(a[16]), .B(n1754), .Z(n74) );
  COND2X1 U1346 ( .A(n77), .B(n1157), .C(n1156), .D(n74), .Z(n878) );
  CENX1 U1347 ( .A(n1560), .B(n505), .Z(n476) );
  CENX1 U1348 ( .A(n484), .B(n486), .Z(n1560) );
  CENXL U1349 ( .A(n1715), .B(b[27]), .Z(n1349) );
  CENXL U1350 ( .A(n1719), .B(b[27]), .Z(n1316) );
  CENXL U1351 ( .A(n1729), .B(b[27]), .Z(n1285) );
  CIVX4 U1352 ( .A(n1739), .Z(n1736) );
  COND2X1 U1353 ( .A(n44), .B(n1245), .C(n1244), .D(n1582), .Z(n962) );
  CENXL U1354 ( .A(n1732), .B(n1392), .Z(n1295) );
  CENXL U1355 ( .A(n1732), .B(n1391), .Z(n1294) );
  CENXL U1356 ( .A(n1732), .B(n1393), .Z(n1296) );
  CENXL U1357 ( .A(n1732), .B(n1394), .Z(n1297) );
  CENXL U1358 ( .A(n1715), .B(b[26]), .Z(n1350) );
  CENXL U1359 ( .A(n1728), .B(b[26]), .Z(n1286) );
  CENXL U1360 ( .A(n1719), .B(b[26]), .Z(n1317) );
  CENX2 U1361 ( .A(n86), .B(a[22]), .Z(n95) );
  CENXL U1362 ( .A(n1729), .B(n1386), .Z(n1289) );
  CENXL U1363 ( .A(n1729), .B(n1388), .Z(n1291) );
  CENXL U1364 ( .A(n1729), .B(n1389), .Z(n1292) );
  CEOX1 U1365 ( .A(a[20]), .B(n86), .Z(n1415) );
  CFA1XL U1366 ( .A(n968), .B(n1076), .CI(n1018), .CO(n727), .S(n728) );
  CNR2IXL U1367 ( .B(n1710), .A(n110), .Z(n824) );
  COND2XL U1368 ( .A(n1096), .B(n112), .C(n110), .D(n1095), .Z(n823) );
  COND2XL U1369 ( .A(n112), .B(n1094), .C(n110), .D(n1093), .Z(n821) );
  CIVX2 U1370 ( .A(n195), .Z(n194) );
  COND2X1 U1371 ( .A(n84), .B(n1145), .C(n1144), .D(n82), .Z(n867) );
  CNIVX1 U1372 ( .A(n962), .Z(n1561) );
  CND2X2 U1373 ( .A(n1412), .B(n105), .Z(n107) );
  CFA1XL U1374 ( .A(n820), .B(n832), .CI(n826), .CO(n409), .S(n410) );
  CENX4 U1375 ( .A(n1763), .B(a[20]), .Z(n89) );
  CIVX4 U1376 ( .A(n1767), .Z(n1763) );
  COND2X1 U1377 ( .A(n53), .B(n1223), .C(n1222), .D(n1583), .Z(n941) );
  CENX2 U1378 ( .A(n1562), .B(n1563), .Z(product[30]) );
  CAN2X2 U1379 ( .A(n1605), .B(n160), .Z(n1562) );
  CANR1X2 U1380 ( .A(n1603), .B(n166), .C(n163), .Z(n1563) );
  CND2X2 U1381 ( .A(n95), .B(n1414), .Z(n97) );
  CIVXL U1382 ( .A(n1676), .Z(n304) );
  CENXL U1383 ( .A(n257), .B(n133), .Z(product[17]) );
  CANR1X1 U1384 ( .A(n182), .B(n169), .C(n170), .Z(n168) );
  CIVX1 U1385 ( .A(n195), .Z(n1569) );
  CNIVX2 U1386 ( .A(n71), .Z(n1590) );
  CNIVX4 U1387 ( .A(n71), .Z(n1686) );
  CIVX1 U1388 ( .A(n71), .Z(n1762) );
  CEOX2 U1389 ( .A(a[6]), .B(n1737), .Z(n1422) );
  CEOX2 U1390 ( .A(n1730), .B(a[6]), .Z(n1608) );
  COND2X1 U1391 ( .A(n1552), .B(n1108), .C(n100), .D(n1107), .Z(n833) );
  CENX4 U1392 ( .A(n1707), .B(a[24]), .Z(n100) );
  CENXL U1393 ( .A(n1730), .B(n1399), .Z(n1302) );
  CENXL U1394 ( .A(n1749), .B(n1399), .Z(n1221) );
  CENXL U1395 ( .A(n1742), .B(n1399), .Z(n1246) );
  CENXL U1396 ( .A(n1716), .B(n1399), .Z(n1366) );
  CENXL U1397 ( .A(n1724), .B(n1399), .Z(n1333) );
  CENXL U1398 ( .A(n86), .B(n1399), .Z(n1126) );
  CENXL U1399 ( .A(n1765), .B(n1399), .Z(n1141) );
  CENXL U1400 ( .A(n1735), .B(n1399), .Z(n1273) );
  CENXL U1401 ( .A(n1754), .B(n1399), .Z(n1177) );
  CIVXL U1402 ( .A(n996), .Z(n1564) );
  CIVX1 U1403 ( .A(n1564), .Z(n1565) );
  CENX2 U1404 ( .A(n166), .B(n121), .Z(product[29]) );
  COND1X1 U1405 ( .A(n179), .B(n171), .C(n172), .Z(n170) );
  CHA1XL U1406 ( .A(n883), .B(n857), .CO(n581), .S(n582) );
  COND2XL U1407 ( .A(n1552), .B(n1106), .C(n100), .D(n1105), .Z(n831) );
  COND2XL U1408 ( .A(n1552), .B(n1107), .C(n100), .D(n1106), .Z(n832) );
  COND2XL U1409 ( .A(n1552), .B(n1110), .C(n100), .D(n1109), .Z(n835) );
  COND2XL U1410 ( .A(n102), .B(n1109), .C(n100), .D(n1108), .Z(n834) );
  CANR1X2 U1411 ( .A(n284), .B(n292), .C(n285), .Z(n283) );
  COND1X1 U1412 ( .A(n290), .B(n1682), .C(n1681), .Z(n285) );
  CNR2X1 U1413 ( .A(n198), .B(n214), .Z(n196) );
  CND2X1 U1414 ( .A(n1604), .B(n347), .Z(n214) );
  CNR2XL U1415 ( .A(n1160), .B(n74), .Z(n1592) );
  CIVX2 U1416 ( .A(n1762), .Z(n1760) );
  CENXL U1417 ( .A(n1715), .B(b[25]), .Z(n1351) );
  CENXL U1418 ( .A(n1728), .B(b[25]), .Z(n1287) );
  CENXL U1419 ( .A(n1736), .B(b[25]), .Z(n1258) );
  CENXL U1420 ( .A(n1720), .B(b[25]), .Z(n1318) );
  CENXL U1421 ( .A(n1764), .B(n1401), .Z(n1143) );
  CENXL U1422 ( .A(n1764), .B(n1402), .Z(n1144) );
  CENXL U1423 ( .A(n1764), .B(n1702), .Z(n1148) );
  CENXL U1424 ( .A(n1764), .B(n1700), .Z(n1149) );
  CIVXL U1425 ( .A(n171), .Z(n340) );
  CNR2X2 U1426 ( .A(n440), .B(n465), .Z(n171) );
  CIVX4 U1427 ( .A(n1727), .Z(n1723) );
  CND2X1 U1428 ( .A(n466), .B(n491), .Z(n179) );
  COND2X1 U1429 ( .A(n77), .B(n1159), .C(n1158), .D(n74), .Z(n880) );
  CENXL U1430 ( .A(n1761), .B(n1399), .Z(n1158) );
  CIVX4 U1431 ( .A(n1759), .Z(n1754) );
  CANR1X1 U1432 ( .A(n265), .B(n246), .C(n247), .Z(n1566) );
  COAN1X1 U1433 ( .A(n233), .B(n1566), .C(n234), .Z(n1567) );
  CIVX4 U1434 ( .A(n63), .Z(n1759) );
  COND2X1 U1435 ( .A(n36), .B(n1269), .C(n1268), .D(n33), .Z(n985) );
  CNR2X2 U1436 ( .A(n660), .B(n675), .Z(n248) );
  CANR1X1 U1437 ( .A(n1601), .B(n244), .C(n241), .Z(n239) );
  CENX2 U1438 ( .A(n1580), .B(n239), .Z(product[20]) );
  COND2XL U1439 ( .A(n97), .B(n1116), .C(n1115), .D(n95), .Z(n840) );
  COND2XL U1440 ( .A(n97), .B(n1119), .C(n1118), .D(n95), .Z(n843) );
  COND2XL U1441 ( .A(n97), .B(n1120), .C(n1119), .D(n95), .Z(n844) );
  COND2XL U1442 ( .A(n97), .B(n1121), .C(n95), .D(n1120), .Z(n845) );
  CNR2IX1 U1443 ( .B(n1710), .A(n95), .Z(n848) );
  CANR1X1 U1444 ( .A(n174), .B(n194), .C(n175), .Z(n173) );
  CNR2IXL U1445 ( .B(n181), .A(n1555), .Z(n174) );
  CNR2X2 U1446 ( .A(n187), .B(n192), .Z(n181) );
  CNR2X2 U1447 ( .A(n516), .B(n539), .Z(n192) );
  CENXL U1448 ( .A(n1715), .B(b[24]), .Z(n1352) );
  CENXL U1449 ( .A(n1728), .B(b[24]), .Z(n1288) );
  CENXL U1450 ( .A(n1720), .B(b[24]), .Z(n1319) );
  CENXL U1451 ( .A(n1734), .B(b[24]), .Z(n1259) );
  CIVX4 U1452 ( .A(n1750), .Z(n1749) );
  CIVX3 U1453 ( .A(n48), .Z(n1750) );
  CND2X2 U1454 ( .A(n1568), .B(n1569), .Z(n1570) );
  CND2X2 U1455 ( .A(n1570), .B(n168), .Z(n166) );
  CIVX2 U1456 ( .A(n167), .Z(n1568) );
  CND2X1 U1457 ( .A(n169), .B(n181), .Z(n167) );
  CANR1X1 U1458 ( .A(n228), .B(n1604), .C(n221), .Z(n215) );
  CIVXL U1459 ( .A(n226), .Z(n228) );
  COND1X1 U1460 ( .A(n215), .B(n198), .C(n199), .Z(n197) );
  CNR2X2 U1461 ( .A(n492), .B(n515), .Z(n187) );
  CEOX2 U1462 ( .A(n123), .B(n180), .Z(product[27]) );
  CENX4 U1463 ( .A(n1736), .B(a[8]), .Z(n1582) );
  CEOX2 U1464 ( .A(n122), .B(n173), .Z(product[28]) );
  COND1X1 U1465 ( .A(n248), .B(n252), .C(n249), .Z(n247) );
  COND2X1 U1466 ( .A(n77), .B(n1167), .C(n1166), .D(n74), .Z(n888) );
  CIVX3 U1467 ( .A(n3), .Z(n1718) );
  COND2X1 U1468 ( .A(n18), .B(n1340), .C(n1339), .D(n15), .Z(n1054) );
  COND2XL U1469 ( .A(n36), .B(n1260), .C(n1259), .D(n33), .Z(n976) );
  COND2XL U1470 ( .A(n36), .B(n1259), .C(n1258), .D(n33), .Z(n975) );
  COND2XL U1471 ( .A(n36), .B(n1279), .C(n1278), .D(n33), .Z(n995) );
  COND2XL U1472 ( .A(n36), .B(n1275), .C(n1274), .D(n33), .Z(n991) );
  COND2XL U1473 ( .A(n36), .B(n1274), .C(n1273), .D(n33), .Z(n990) );
  COND2XL U1474 ( .A(n36), .B(n1262), .C(n1261), .D(n33), .Z(n978) );
  COND2XL U1475 ( .A(n36), .B(n1261), .C(n1260), .D(n33), .Z(n977) );
  COND2XL U1476 ( .A(n36), .B(n1282), .C(n1281), .D(n33), .Z(n998) );
  COND2XL U1477 ( .A(n36), .B(n1273), .C(n1272), .D(n33), .Z(n989) );
  COND2XL U1478 ( .A(n36), .B(n1272), .C(n1271), .D(n33), .Z(n988) );
  COND2XL U1479 ( .A(n36), .B(n1270), .C(n1269), .D(n33), .Z(n986) );
  COND2XL U1480 ( .A(n36), .B(n1271), .C(n1270), .D(n33), .Z(n987) );
  COND2XL U1481 ( .A(n36), .B(n1277), .C(n1276), .D(n33), .Z(n993) );
  COND2XL U1482 ( .A(n36), .B(n1264), .C(n1263), .D(n33), .Z(n980) );
  COND2XL U1483 ( .A(n36), .B(n1281), .C(n1280), .D(n33), .Z(n997) );
  COND2XL U1484 ( .A(n36), .B(n1276), .C(n1275), .D(n33), .Z(n992) );
  COND2XL U1485 ( .A(n1283), .B(n36), .C(n1282), .D(n33), .Z(n999) );
  COND2XL U1486 ( .A(n36), .B(n1263), .C(n1262), .D(n33), .Z(n979) );
  COND2XL U1487 ( .A(n36), .B(n1267), .C(n1266), .D(n33), .Z(n983) );
  COND2XL U1488 ( .A(n36), .B(n1278), .C(n1277), .D(n33), .Z(n994) );
  COND2XL U1489 ( .A(n36), .B(n1280), .C(n1279), .D(n33), .Z(n996) );
  CND2X1 U1490 ( .A(n504), .B(n525), .Z(n1571) );
  CND2X1 U1491 ( .A(n504), .B(n527), .Z(n1572) );
  CND2X1 U1492 ( .A(n525), .B(n527), .Z(n1573) );
  CND3X1 U1493 ( .A(n1571), .B(n1572), .C(n1573), .Z(n497) );
  CIVX2 U1494 ( .A(n1753), .Z(n1752) );
  CIVX1 U1495 ( .A(n265), .Z(n264) );
  CANR1X1 U1496 ( .A(n343), .B(n194), .C(n191), .Z(n189) );
  CHA1XL U1497 ( .A(n927), .B(n812), .CO(n741), .S(n742) );
  CFA1X1 U1498 ( .A(n807), .B(n959), .CI(n899), .CO(n579), .S(n580) );
  CENXL U1499 ( .A(n1717), .B(n1396), .Z(n1363) );
  CENXL U1500 ( .A(n1717), .B(n1393), .Z(n1360) );
  CENXL U1501 ( .A(n1717), .B(n1395), .Z(n1362) );
  CENXL U1502 ( .A(n1717), .B(n1394), .Z(n1361) );
  CND2IXL U1503 ( .B(n1710), .A(n1717), .Z(n1377) );
  CENXL U1504 ( .A(n1709), .B(n1717), .Z(n1376) );
  CENXL U1505 ( .A(n1717), .B(n1392), .Z(n1359) );
  CENXL U1506 ( .A(n1717), .B(n1397), .Z(n1364) );
  CENX4 U1507 ( .A(n1741), .B(a[10]), .Z(n1583) );
  COND2X1 U1508 ( .A(n53), .B(n1218), .C(n1217), .D(n1583), .Z(n936) );
  COND2X1 U1509 ( .A(n53), .B(n1216), .C(n1215), .D(n1583), .Z(n934) );
  COND2X1 U1510 ( .A(n53), .B(n1230), .C(n1229), .D(n1583), .Z(n948) );
  CENX4 U1511 ( .A(n1723), .B(a[4]), .Z(n24) );
  COND2X1 U1512 ( .A(n27), .B(n1292), .C(n1291), .D(n24), .Z(n1007) );
  COND2X1 U1513 ( .A(n61), .B(n1202), .C(n1201), .D(n1550), .Z(n921) );
  CND2X4 U1514 ( .A(n1419), .B(n58), .Z(n61) );
  CENXL U1515 ( .A(n204), .B(n126), .Z(product[24]) );
  CENXL U1516 ( .A(n1760), .B(n1401), .Z(n1160) );
  CENXL U1517 ( .A(n1763), .B(n1403), .Z(n1145) );
  CENX2 U1518 ( .A(n213), .B(n127), .Z(product[23]) );
  COND1X1 U1519 ( .A(n214), .B(n1567), .C(n215), .Z(n213) );
  CENXL U1520 ( .A(n1720), .B(n1387), .Z(n1321) );
  COND2X1 U1521 ( .A(n97), .B(n1122), .C(n95), .D(n1121), .Z(n846) );
  COND2X1 U1522 ( .A(n69), .B(n1178), .C(n1177), .D(n66), .Z(n898) );
  COND2X1 U1523 ( .A(n69), .B(n1179), .C(n1178), .D(n66), .Z(n899) );
  COND2X1 U1524 ( .A(n69), .B(n1173), .C(n1172), .D(n66), .Z(n893) );
  CENXL U1525 ( .A(n1743), .B(n1395), .Z(n1242) );
  CENXL U1526 ( .A(n1743), .B(n1394), .Z(n1241) );
  CENXL U1527 ( .A(n1743), .B(n1393), .Z(n1240) );
  CENXL U1528 ( .A(n1743), .B(n1392), .Z(n1239) );
  CNIVX2 U1529 ( .A(n1008), .Z(n1574) );
  COND2X1 U1530 ( .A(n27), .B(n1290), .C(n1289), .D(n24), .Z(n1005) );
  CENXL U1531 ( .A(n1729), .B(n1387), .Z(n1290) );
  CEOX2 U1532 ( .A(a[12]), .B(n1752), .Z(n1419) );
  CENXL U1533 ( .A(n1752), .B(n1396), .Z(n1195) );
  CENXL U1534 ( .A(n1752), .B(n1395), .Z(n1194) );
  CENXL U1535 ( .A(n1752), .B(n1394), .Z(n1193) );
  CENXL U1536 ( .A(n1710), .B(n1752), .Z(n1208) );
  CND2IXL U1537 ( .B(n1710), .A(n1752), .Z(n1209) );
  CENXL U1538 ( .A(n1752), .B(n1392), .Z(n1191) );
  CENXL U1539 ( .A(n1752), .B(n1393), .Z(n1192) );
  CENXL U1540 ( .A(n1752), .B(n1391), .Z(n1190) );
  CFA1X1 U1541 ( .A(n881), .B(n1007), .CI(n915), .CO(n533), .S(n534) );
  CND2X2 U1542 ( .A(n516), .B(n539), .Z(n193) );
  CFA1X1 U1543 ( .A(n868), .B(n982), .CI(n898), .CO(n557), .S(n558) );
  COND1X1 U1544 ( .A(n1555), .B(n184), .C(n179), .Z(n175) );
  CIVX8 U1545 ( .A(n1718), .Z(n1716) );
  CFA1XL U1546 ( .A(n992), .B(n741), .CI(n1046), .CO(n725), .S(n726) );
  CFA1XL U1547 ( .A(n1000), .B(n1054), .CI(n1026), .CO(n793), .S(n794) );
  CFA1XL U1548 ( .A(n1025), .B(n1083), .CI(n1053), .CO(n787), .S(n788) );
  CIVX4 U1549 ( .A(n1753), .Z(n1751) );
  CENXL U1550 ( .A(n1751), .B(n1397), .Z(n1196) );
  CENXL U1551 ( .A(n1751), .B(n1401), .Z(n1200) );
  CENXL U1552 ( .A(n1751), .B(n1402), .Z(n1201) );
  CENXL U1553 ( .A(n1751), .B(n1398), .Z(n1197) );
  CENXL U1554 ( .A(n1751), .B(n1403), .Z(n1202) );
  CENXL U1555 ( .A(n1751), .B(n1399), .Z(n1198) );
  CENXL U1556 ( .A(n1751), .B(n1711), .Z(n1207) );
  CANR1X2 U1557 ( .A(n196), .B(n232), .C(n197), .Z(n195) );
  CENX4 U1558 ( .A(n1751), .B(a[14]), .Z(n66) );
  CIVX4 U1559 ( .A(n1750), .Z(n1748) );
  CND2X2 U1560 ( .A(n89), .B(n1415), .Z(n91) );
  CND2XL U1561 ( .A(n802), .B(n1057), .Z(n328) );
  CND2X1 U1562 ( .A(n1575), .B(n1576), .Z(n807) );
  COR2XL U1563 ( .A(n1439), .B(n97), .Z(n1576) );
  CIVX4 U1564 ( .A(n1701), .Z(n1702) );
  COND1XL U1565 ( .A(n329), .B(n327), .C(n328), .Z(n326) );
  COND1XL U1566 ( .A(n321), .B(n319), .C(n320), .Z(n318) );
  CND2IX1 U1567 ( .B(n311), .A(n312), .Z(n143) );
  COND1X1 U1568 ( .A(n233), .B(n245), .C(n234), .Z(n232) );
  CND2X1 U1569 ( .A(n1603), .B(n165), .Z(n121) );
  COR2X1 U1570 ( .A(n562), .B(n583), .Z(n1602) );
  COR2X1 U1571 ( .A(n1591), .B(n1592), .Z(n882) );
  CNR2X1 U1572 ( .A(n77), .B(n1161), .Z(n1591) );
  CIVX2 U1573 ( .A(n1714), .Z(n1586) );
  CENX1 U1574 ( .A(a[18]), .B(n1766), .Z(n1581) );
  CIVX4 U1575 ( .A(n1703), .Z(n1704) );
  COR2XL U1576 ( .A(n1124), .B(n95), .Z(n1575) );
  CND2IXL U1577 ( .B(n1710), .A(n1707), .Z(n1124) );
  CIVXL U1578 ( .A(n1707), .Z(n1439) );
  COND1X1 U1579 ( .A(n311), .B(n313), .C(n312), .Z(n310) );
  CANR1X1 U1580 ( .A(n326), .B(n1597), .C(n323), .Z(n321) );
  CANR1X1 U1581 ( .A(n318), .B(n1596), .C(n315), .Z(n313) );
  CND2XL U1582 ( .A(n1596), .B(n317), .Z(n144) );
  CND2XL U1583 ( .A(n1598), .B(n333), .Z(n148) );
  CNR2XL U1584 ( .A(n744), .B(n753), .Z(n286) );
  CND2XL U1585 ( .A(n764), .B(n771), .Z(n298) );
  CND2XL U1586 ( .A(n772), .B(n779), .Z(n303) );
  CND2IXL U1587 ( .B(n319), .A(n320), .Z(n145) );
  CND2IXL U1588 ( .B(n327), .A(n328), .Z(n147) );
  CENX1 U1589 ( .A(n1577), .B(n264), .Z(product[16]) );
  CAN2XL U1590 ( .A(n352), .B(n259), .Z(n1577) );
  CENX1 U1591 ( .A(n1578), .B(n1567), .Z(product[21]) );
  CAN2XL U1592 ( .A(n347), .B(n226), .Z(n1578) );
  CANR1X1 U1593 ( .A(n246), .B(n265), .C(n247), .Z(n245) );
  CANR1X1 U1594 ( .A(n261), .B(n1599), .C(n254), .Z(n252) );
  CIVX1 U1595 ( .A(n256), .Z(n254) );
  CND2XL U1596 ( .A(n1600), .B(n1601), .Z(n233) );
  CND3X1 U1597 ( .A(n1690), .B(n1691), .C(n1692), .Z(n475) );
  CND2XL U1598 ( .A(n1599), .B(n256), .Z(n133) );
  CND2XL U1599 ( .A(n1601), .B(n243), .Z(n131) );
  CND2XL U1600 ( .A(n1604), .B(n223), .Z(n128) );
  CIVXL U1601 ( .A(n223), .Z(n221) );
  CND2XL U1602 ( .A(n343), .B(n193), .Z(n125) );
  CND2XL U1603 ( .A(n344), .B(n203), .Z(n126) );
  CENX1 U1604 ( .A(n1579), .B(n189), .Z(product[26]) );
  CAN2XL U1605 ( .A(n342), .B(n188), .Z(n1579) );
  CAN2XL U1606 ( .A(n1600), .B(n238), .Z(n1580) );
  CND2XL U1607 ( .A(n350), .B(n249), .Z(n132) );
  CIVXL U1608 ( .A(n215), .Z(n217) );
  CND2XL U1609 ( .A(n1599), .B(n352), .Z(n251) );
  COR2XL U1610 ( .A(n1088), .B(n1058), .Z(n1598) );
  CND2IXL U1611 ( .B(n335), .A(n336), .Z(n149) );
  CANR1X1 U1612 ( .A(n1607), .B(n274), .C(n269), .Z(n267) );
  COND1X1 U1613 ( .A(n283), .B(n266), .C(n267), .Z(n265) );
  CND2XL U1614 ( .A(n273), .B(n1607), .Z(n266) );
  CNR2IXL U1615 ( .B(n1710), .A(n89), .Z(n860) );
  CNR2IXL U1616 ( .B(n1710), .A(n82), .Z(n874) );
  CNR2IXL U1617 ( .B(n1710), .A(n66), .Z(n908) );
  CND2X1 U1618 ( .A(n562), .B(n583), .Z(n212) );
  CEOXL U1619 ( .A(n135), .B(n272), .Z(product[15]) );
  CND2XL U1620 ( .A(n1607), .B(n271), .Z(n135) );
  CEOXL U1621 ( .A(n136), .B(n277), .Z(product[14]) );
  CND2XL U1622 ( .A(n357), .B(n290), .Z(n139) );
  CEOXL U1623 ( .A(n139), .B(n291), .Z(product[11]) );
  CNR2IXL U1624 ( .B(n1710), .A(n15), .Z(n1058) );
  CNR2XL U1625 ( .A(n275), .B(n280), .Z(n273) );
  CND2XL U1626 ( .A(n355), .B(n281), .Z(n137) );
  CNR2IXL U1627 ( .B(n1710), .A(n114), .Z(n820) );
  CNR2IXL U1628 ( .B(n1710), .A(n33), .Z(n1000) );
  CNR2IXL U1629 ( .B(n1710), .A(n1713), .Z(product[0]) );
  CENX4 U1630 ( .A(n1686), .B(a[18]), .Z(n82) );
  CND2IX4 U1631 ( .B(n1581), .A(n82), .Z(n84) );
  CENX4 U1632 ( .A(n1716), .B(a[2]), .Z(n15) );
  CNIVX2 U1633 ( .A(n116), .Z(n1709) );
  CIVX3 U1634 ( .A(n1608), .Z(n33) );
  CND2IX4 U1635 ( .B(n1611), .A(n1583), .Z(n53) );
  CND2X4 U1636 ( .A(n1424), .B(n15), .Z(n18) );
  CEOX2 U1637 ( .A(a[2]), .B(n1723), .Z(n1424) );
  CENXL U1638 ( .A(a[8]), .B(n1744), .Z(n1584) );
  CNR2X2 U1639 ( .A(n1587), .B(n1586), .Z(n1585) );
  CANR1X1 U1640 ( .A(n301), .B(n1684), .C(n296), .Z(n294) );
  CIVX3 U1641 ( .A(n1699), .Z(n1700) );
  CND2IX4 U1642 ( .B(n1588), .A(n66), .Z(n69) );
  CND2IX4 U1643 ( .B(n1589), .A(n24), .Z(n27) );
  CENXL U1644 ( .A(a[4]), .B(n21), .Z(n1589) );
  CIVX2 U1645 ( .A(n79), .Z(n1767) );
  CND2XL U1646 ( .A(n1618), .B(n1616), .Z(n276) );
  CIVX2 U1647 ( .A(n55), .Z(n1753) );
  CIVX3 U1648 ( .A(n1705), .Z(n1706) );
  CENX1 U1649 ( .A(n1761), .B(n1402), .Z(n1161) );
  CENX1 U1650 ( .A(n142), .B(n310), .Z(product[8]) );
  CND2X1 U1651 ( .A(n1593), .B(n309), .Z(n142) );
  CANR1XL U1652 ( .A(n1593), .B(n310), .C(n307), .Z(n305) );
  CANR1XL U1653 ( .A(n334), .B(n1598), .C(n331), .Z(n329) );
  CENX1 U1654 ( .A(n144), .B(n318), .Z(product[6]) );
  CENX1 U1655 ( .A(n148), .B(n334), .Z(product[2]) );
  CENX1 U1656 ( .A(n146), .B(n326), .Z(product[4]) );
  CND2X1 U1657 ( .A(n1597), .B(n325), .Z(n146) );
  CND2X1 U1658 ( .A(n780), .B(n785), .Z(n309) );
  COR2X1 U1659 ( .A(n780), .B(n785), .Z(n1593) );
  CND2XL U1660 ( .A(n744), .B(n753), .Z(n287) );
  COR2X1 U1661 ( .A(n764), .B(n771), .Z(n1594) );
  COR2X1 U1662 ( .A(n772), .B(n779), .Z(n1595) );
  CND2X1 U1663 ( .A(n1602), .B(n212), .Z(n127) );
  CANR1X1 U1664 ( .A(n241), .B(n1600), .C(n236), .Z(n234) );
  CENX1 U1665 ( .A(n194), .B(n125), .Z(product[25]) );
  CND2X1 U1666 ( .A(n1554), .B(n179), .Z(n123) );
  COND1XL U1667 ( .A(n258), .B(n264), .C(n259), .Z(n257) );
  CENX1 U1668 ( .A(n244), .B(n131), .Z(product[19]) );
  CND2X1 U1669 ( .A(n216), .B(n1602), .Z(n205) );
  CANR1XL U1670 ( .A(n1602), .B(n217), .C(n210), .Z(n206) );
  CANR1XL U1671 ( .A(n1556), .B(n166), .C(n154), .Z(n152) );
  CNR2X1 U1672 ( .A(n786), .B(n791), .Z(n311) );
  CNR2X1 U1673 ( .A(n796), .B(n799), .Z(n319) );
  CANR1XL U1674 ( .A(n163), .B(n1605), .C(n158), .Z(n156) );
  CNR2X1 U1675 ( .A(n802), .B(n1057), .Z(n327) );
  CND2X1 U1676 ( .A(n786), .B(n791), .Z(n312) );
  CND2X1 U1677 ( .A(n796), .B(n799), .Z(n320) );
  CND2X1 U1678 ( .A(n792), .B(n795), .Z(n317) );
  CND2X1 U1679 ( .A(n1089), .B(n818), .Z(n336) );
  CND2X1 U1680 ( .A(n800), .B(n801), .Z(n325) );
  CND2X1 U1681 ( .A(n1088), .B(n1058), .Z(n333) );
  COR2X1 U1682 ( .A(n792), .B(n795), .Z(n1596) );
  COR2X1 U1683 ( .A(n800), .B(n801), .Z(n1597) );
  CNR2XL U1684 ( .A(n1089), .B(n818), .Z(n335) );
  COND1XL U1685 ( .A(n281), .B(n275), .C(n276), .Z(n274) );
  CNR2X1 U1686 ( .A(n692), .B(n705), .Z(n258) );
  COR2X1 U1687 ( .A(n676), .B(n691), .Z(n1599) );
  COR2X1 U1688 ( .A(n624), .B(n641), .Z(n1600) );
  COR2X1 U1689 ( .A(n642), .B(n659), .Z(n1601) );
  CND2X1 U1690 ( .A(n692), .B(n705), .Z(n259) );
  CND2X1 U1691 ( .A(n660), .B(n675), .Z(n249) );
  CND2X1 U1692 ( .A(n642), .B(n659), .Z(n243) );
  CND2X1 U1693 ( .A(n624), .B(n641), .Z(n238) );
  CND2X1 U1694 ( .A(n676), .B(n691), .Z(n256) );
  CENX1 U1695 ( .A(n1709), .B(n1726), .Z(n1343) );
  COND2X1 U1696 ( .A(n84), .B(n1143), .C(n1142), .D(n82), .Z(n865) );
  CENX1 U1697 ( .A(n1736), .B(n1711), .Z(n1282) );
  CENX1 U1698 ( .A(n1748), .B(n1706), .Z(n1226) );
  CENX1 U1699 ( .A(n86), .B(n1704), .Z(n1132) );
  CENX1 U1700 ( .A(n1758), .B(n1704), .Z(n1183) );
  CENX1 U1701 ( .A(n1756), .B(n1706), .Z(n1182) );
  CENX1 U1702 ( .A(n1716), .B(n1706), .Z(n1371) );
  CENX1 U1703 ( .A(n1716), .B(n1700), .Z(n1374) );
  CENX1 U1704 ( .A(n1716), .B(n1704), .Z(n1372) );
  CENX1 U1705 ( .A(n1716), .B(n1702), .Z(n1373) );
  CENX1 U1706 ( .A(n1716), .B(n1712), .Z(n1375) );
  CND2X1 U1707 ( .A(n354), .B(n276), .Z(n136) );
  CANR1XL U1708 ( .A(n355), .B(n282), .C(n279), .Z(n277) );
  CANR1XL U1709 ( .A(n273), .B(n282), .C(n274), .Z(n272) );
  CENX1 U1710 ( .A(n1741), .B(n1700), .Z(n1254) );
  CENX1 U1711 ( .A(n1757), .B(n1700), .Z(n1185) );
  CENX1 U1712 ( .A(n1741), .B(n1711), .Z(n1255) );
  CENX1 U1713 ( .A(n1757), .B(n1711), .Z(n1186) );
  CENX1 U1714 ( .A(n1723), .B(n1712), .Z(n1342) );
  CENX1 U1715 ( .A(n1758), .B(n1702), .Z(n1184) );
  CENX1 U1716 ( .A(n282), .B(n137), .Z(product[13]) );
  CENX1 U1717 ( .A(n1709), .B(n86), .Z(n1136) );
  CIVX2 U1718 ( .A(n1733), .Z(n1729) );
  CENX1 U1719 ( .A(n1741), .B(n1702), .Z(n1253) );
  CIVX2 U1720 ( .A(n1718), .Z(n1715) );
  CENX1 U1721 ( .A(n1735), .B(n1704), .Z(n1279) );
  CENX1 U1722 ( .A(n86), .B(n1706), .Z(n1131) );
  CENX1 U1723 ( .A(n1704), .B(n1707), .Z(n1119) );
  CENX1 U1724 ( .A(n1735), .B(n1702), .Z(n1280) );
  CENX1 U1725 ( .A(n1735), .B(n1700), .Z(n1281) );
  CENX1 U1726 ( .A(n1763), .B(n1706), .Z(n1146) );
  CENX1 U1727 ( .A(n1700), .B(n86), .Z(n1134) );
  CENX1 U1728 ( .A(n1763), .B(n1704), .Z(n1147) );
  CENX1 U1729 ( .A(n1702), .B(n86), .Z(n1133) );
  CENX1 U1730 ( .A(n1735), .B(n1706), .Z(n1278) );
  CENX1 U1731 ( .A(n1686), .B(n1706), .Z(n1163) );
  CIVX2 U1732 ( .A(n1745), .Z(n1740) );
  CENX1 U1733 ( .A(n1711), .B(n86), .Z(n1135) );
  CENX1 U1734 ( .A(n1702), .B(n1707), .Z(n1120) );
  CENX1 U1735 ( .A(n1706), .B(n1708), .Z(n1107) );
  CENX1 U1736 ( .A(n1700), .B(n1708), .Z(n1110) );
  CENX1 U1737 ( .A(n1711), .B(n1708), .Z(n1111) );
  CENX1 U1738 ( .A(n1700), .B(n1707), .Z(n1121) );
  CENX1 U1739 ( .A(n1704), .B(n1708), .Z(n1108) );
  CENX1 U1740 ( .A(n1702), .B(n1708), .Z(n1109) );
  CENX1 U1741 ( .A(n1706), .B(n1707), .Z(n1118) );
  CENX1 U1742 ( .A(n1748), .B(n1704), .Z(n1227) );
  CENX1 U1743 ( .A(n1686), .B(n1704), .Z(n1164) );
  CENX1 U1744 ( .A(n1711), .B(n1707), .Z(n1122) );
  CENX1 U1745 ( .A(n1710), .B(n1729), .Z(n1312) );
  CENX1 U1746 ( .A(n1709), .B(n1749), .Z(n1231) );
  CENX1 U1747 ( .A(n1709), .B(n1708), .Z(n1112) );
  CENX1 U1748 ( .A(n1729), .B(n1712), .Z(n1311) );
  CENX1 U1749 ( .A(n1751), .B(n1700), .Z(n1206) );
  CENX1 U1750 ( .A(n1751), .B(n1702), .Z(n1205) );
  CENX1 U1751 ( .A(n1751), .B(n1704), .Z(n1204) );
  CENX1 U1752 ( .A(n1729), .B(n1706), .Z(n1307) );
  CENX1 U1753 ( .A(n1729), .B(n1704), .Z(n1308) );
  CENX1 U1754 ( .A(n1760), .B(n1700), .Z(n1166) );
  CENX1 U1755 ( .A(n1740), .B(n1704), .Z(n1252) );
  CENX1 U1756 ( .A(n1711), .B(n1761), .Z(n1167) );
  CENX1 U1757 ( .A(n1742), .B(n1706), .Z(n1251) );
  CENX1 U1758 ( .A(n1729), .B(n1700), .Z(n1310) );
  CENX1 U1759 ( .A(n1748), .B(n1700), .Z(n1229) );
  CENX1 U1760 ( .A(n1760), .B(n1702), .Z(n1165) );
  CENX1 U1761 ( .A(n1729), .B(n1702), .Z(n1309) );
  CENX1 U1762 ( .A(n1748), .B(n1702), .Z(n1228) );
  CENX1 U1763 ( .A(n1748), .B(n1711), .Z(n1230) );
  CENX1 U1764 ( .A(n1751), .B(n1706), .Z(n1203) );
  CNR2X1 U1765 ( .A(n604), .B(n623), .Z(n225) );
  CENX1 U1766 ( .A(n1709), .B(n1707), .Z(n1123) );
  CIVX2 U1767 ( .A(n1718), .Z(n1717) );
  CENX1 U1768 ( .A(n1710), .B(n1761), .Z(n1168) );
  COND2X1 U1769 ( .A(n36), .B(n1268), .C(n1267), .D(n33), .Z(n984) );
  COR2X1 U1770 ( .A(n412), .B(n439), .Z(n1603) );
  CNR2X1 U1771 ( .A(n540), .B(n561), .Z(n202) );
  CND2X1 U1772 ( .A(n604), .B(n623), .Z(n226) );
  COR2X1 U1773 ( .A(n584), .B(n603), .Z(n1604) );
  COR2X1 U1774 ( .A(n384), .B(n411), .Z(n1605) );
  CND2X1 U1775 ( .A(n492), .B(n515), .Z(n188) );
  CENX1 U1776 ( .A(n1709), .B(n1737), .Z(n1283) );
  CNR2IX1 U1777 ( .B(n1710), .A(n1583), .Z(n950) );
  CND2X1 U1778 ( .A(n584), .B(n603), .Z(n223) );
  CND2X1 U1779 ( .A(n412), .B(n439), .Z(n165) );
  CND2X1 U1780 ( .A(n384), .B(n411), .Z(n160) );
  CND2X1 U1781 ( .A(n540), .B(n561), .Z(n203) );
  CIVX2 U1782 ( .A(n1733), .Z(n1730) );
  COR2X1 U1783 ( .A(n150), .B(n1606), .Z(n119) );
  CAN2X1 U1784 ( .A(n383), .B(n368), .Z(n1606) );
  CNR2X1 U1785 ( .A(n383), .B(n368), .Z(n150) );
  CNR2XL U1786 ( .A(n1682), .B(n289), .Z(n284) );
  CNR2X1 U1787 ( .A(n1613), .B(n1612), .Z(n289) );
  COND1X1 U1788 ( .A(n1676), .B(n293), .C(n294), .Z(n292) );
  CND2XL U1789 ( .A(n1684), .B(n1683), .Z(n293) );
  CNR2X1 U1790 ( .A(n1618), .B(n1616), .Z(n275) );
  COR2X1 U1791 ( .A(n706), .B(n1619), .Z(n1607) );
  CND2X1 U1792 ( .A(n1615), .B(n1614), .Z(n281) );
  CND2X1 U1793 ( .A(n1613), .B(n1612), .Z(n290) );
  CND2X1 U1794 ( .A(n706), .B(n1619), .Z(n271) );
  CENX1 U1795 ( .A(n1735), .B(n1394), .Z(n1268) );
  CENX1 U1796 ( .A(n1735), .B(n1393), .Z(n1267) );
  CENX1 U1797 ( .A(n1752), .B(n1390), .Z(n1189) );
  CENX1 U1798 ( .A(n1725), .B(n1396), .Z(n1330) );
  CENX1 U1799 ( .A(n1725), .B(n1394), .Z(n1328) );
  CENX1 U1800 ( .A(n1735), .B(n1397), .Z(n1271) );
  CENX1 U1801 ( .A(n1735), .B(n1396), .Z(n1270) );
  CENX1 U1802 ( .A(n86), .B(n1402), .Z(n1129) );
  CENX1 U1803 ( .A(n86), .B(n1401), .Z(n1128) );
  CENX1 U1804 ( .A(n1734), .B(n1387), .Z(n1261) );
  CENX1 U1805 ( .A(n1765), .B(n1397), .Z(n1139) );
  CENX1 U1806 ( .A(n1734), .B(n1402), .Z(n1276) );
  CENX1 U1807 ( .A(n1736), .B(n1401), .Z(n1275) );
  CENX1 U1808 ( .A(n1734), .B(n1386), .Z(n1260) );
  CENX1 U1809 ( .A(n1758), .B(n1401), .Z(n1179) );
  CENX1 U1810 ( .A(n1734), .B(n1390), .Z(n1264) );
  CENX1 U1811 ( .A(n1756), .B(n1402), .Z(n1180) );
  CENX1 U1812 ( .A(n1758), .B(n1397), .Z(n1175) );
  CENX1 U1813 ( .A(n86), .B(n1403), .Z(n1130) );
  CENX1 U1814 ( .A(n1755), .B(n1403), .Z(n1181) );
  CENX1 U1815 ( .A(n1735), .B(n1403), .Z(n1277) );
  CENX1 U1816 ( .A(n1735), .B(n1395), .Z(n1269) );
  CENX1 U1817 ( .A(n1716), .B(n1403), .Z(n1370) );
  CENX1 U1818 ( .A(n1715), .B(n1402), .Z(n1369) );
  CENX1 U1819 ( .A(n1403), .B(n1708), .Z(n1106) );
  CENX1 U1820 ( .A(n1716), .B(n1401), .Z(n1368) );
  CENX1 U1821 ( .A(n1716), .B(n1391), .Z(n1358) );
  CENX1 U1822 ( .A(n104), .B(a[28]), .Z(n110) );
  CENX1 U1823 ( .A(n288), .B(n138), .Z(product[12]) );
  CND2XL U1824 ( .A(n356), .B(n1681), .Z(n138) );
  COND1XL U1825 ( .A(n289), .B(n291), .C(n290), .Z(n288) );
  CENX1 U1826 ( .A(n1729), .B(n1402), .Z(n1305) );
  CENX1 U1827 ( .A(n1748), .B(n1403), .Z(n1225) );
  CENX1 U1828 ( .A(n1707), .B(n1401), .Z(n1115) );
  CENX1 U1829 ( .A(n1757), .B(n1400), .Z(n1178) );
  CENX1 U1830 ( .A(n1749), .B(n1394), .Z(n1216) );
  CENX1 U1831 ( .A(n1686), .B(n1403), .Z(n1162) );
  CENX1 U1832 ( .A(n1726), .B(n1393), .Z(n1327) );
  CENX1 U1833 ( .A(n1757), .B(n1396), .Z(n1174) );
  CENX1 U1834 ( .A(n1720), .B(n1386), .Z(n1320) );
  CENX1 U1835 ( .A(n1740), .B(n1401), .Z(n1248) );
  CENX1 U1836 ( .A(n1732), .B(n1403), .Z(n1306) );
  CENX1 U1837 ( .A(n1402), .B(n1707), .Z(n1116) );
  CENX1 U1838 ( .A(n1740), .B(n1397), .Z(n1244) );
  CENX1 U1839 ( .A(n1724), .B(n1400), .Z(n1334) );
  CENX1 U1840 ( .A(n1740), .B(n1402), .Z(n1249) );
  CENX1 U1841 ( .A(n1725), .B(n1397), .Z(n1331) );
  CENX1 U1842 ( .A(n1723), .B(n1392), .Z(n1326) );
  CENX1 U1843 ( .A(n1719), .B(n1390), .Z(n1324) );
  CENX1 U1844 ( .A(n109), .B(a[30]), .Z(n114) );
  CENX1 U1845 ( .A(n1590), .B(n1394), .Z(n1153) );
  CENX1 U1846 ( .A(n141), .B(n304), .Z(product[9]) );
  CND2XL U1847 ( .A(n1683), .B(n1679), .Z(n141) );
  CENX1 U1848 ( .A(n86), .B(n1398), .Z(n1125) );
  CEOX1 U1849 ( .A(n299), .B(n140), .Z(product[10]) );
  CND2XL U1850 ( .A(n1684), .B(n1680), .Z(n140) );
  CANR1XL U1851 ( .A(n1683), .B(n304), .C(n301), .Z(n299) );
  CENX1 U1852 ( .A(n1402), .B(n1708), .Z(n1105) );
  CENX1 U1853 ( .A(n1716), .B(b[31]), .Z(n1345) );
  CENX1 U1854 ( .A(n1609), .B(n1642), .Z(n584) );
  CENX1 U1855 ( .A(n1641), .B(n1640), .Z(n1609) );
  CENX1 U1856 ( .A(n1610), .B(n1639), .Z(n604) );
  CENX1 U1857 ( .A(n1638), .B(n1637), .Z(n1610) );
  CENX1 U1858 ( .A(n1721), .B(n1403), .Z(n1337) );
  CENX1 U1859 ( .A(n1730), .B(n1401), .Z(n1304) );
  CENX1 U1860 ( .A(n1731), .B(n1398), .Z(n1301) );
  CENX1 U1861 ( .A(n1748), .B(n1402), .Z(n1224) );
  CENX1 U1862 ( .A(n1590), .B(n1395), .Z(n1154) );
  CENX1 U1863 ( .A(n1730), .B(n1400), .Z(n1303) );
  CENX1 U1864 ( .A(n1731), .B(n1397), .Z(n1300) );
  CENX1 U1865 ( .A(n1742), .B(n1403), .Z(n1250) );
  CENX1 U1866 ( .A(n1721), .B(n1402), .Z(n1336) );
  CENX1 U1867 ( .A(n1731), .B(n1395), .Z(n1298) );
  CENX1 U1868 ( .A(n1749), .B(n1393), .Z(n1215) );
  CENX1 U1869 ( .A(n1728), .B(n1390), .Z(n1293) );
  CENX1 U1870 ( .A(n1749), .B(n1392), .Z(n1214) );
  CENX1 U1871 ( .A(n1724), .B(n1401), .Z(n1335) );
  CENX1 U1872 ( .A(n1403), .B(n1707), .Z(n1117) );
  CENX1 U1873 ( .A(n1590), .B(n1396), .Z(n1155) );
  CENX1 U1874 ( .A(n1761), .B(n1397), .Z(n1156) );
  CENX1 U1875 ( .A(n1749), .B(n1400), .Z(n1222) );
  CENX1 U1876 ( .A(n1749), .B(n1391), .Z(n1213) );
  CENX1 U1877 ( .A(n1742), .B(n1398), .Z(n1245) );
  CENX1 U1878 ( .A(n1748), .B(n1401), .Z(n1223) );
  CENX1 U1879 ( .A(n1731), .B(n1396), .Z(n1299) );
  CENX1 U1880 ( .A(n1719), .B(b[28]), .Z(n1315) );
  CENX1 U1881 ( .A(n1734), .B(n1389), .Z(n1263) );
  CENX1 U1882 ( .A(n1735), .B(n1388), .Z(n1262) );
  CENX1 U1883 ( .A(n1721), .B(n1389), .Z(n1323) );
  CENX1 U1884 ( .A(n1737), .B(n1392), .Z(n1266) );
  CENX1 U1885 ( .A(n1737), .B(n1391), .Z(n1265) );
  CENX1 U1886 ( .A(n1721), .B(n1388), .Z(n1322) );
  CENX1 U1887 ( .A(n1742), .B(n1391), .Z(n1238) );
  CENX1 U1888 ( .A(n1715), .B(n1390), .Z(n1357) );
  CENX1 U1889 ( .A(n1715), .B(n1389), .Z(n1356) );
  CENX1 U1890 ( .A(n1715), .B(n1388), .Z(n1355) );
  CENX1 U1891 ( .A(n1715), .B(n1387), .Z(n1354) );
  CENX1 U1892 ( .A(n1715), .B(n1386), .Z(n1353) );
  CENX1 U1893 ( .A(n1704), .B(n104), .Z(n1099) );
  CENX1 U1894 ( .A(n1702), .B(n104), .Z(n1100) );
  CENX1 U1895 ( .A(n1700), .B(n109), .Z(n1094) );
  CENX1 U1896 ( .A(n1715), .B(b[29]), .Z(n1347) );
  CENX1 U1897 ( .A(n1711), .B(n104), .Z(n1102) );
  CENX1 U1898 ( .A(n1700), .B(n104), .Z(n1101) );
  CENX1 U1899 ( .A(n1715), .B(b[28]), .Z(n1348) );
  CENX1 U1900 ( .A(n1715), .B(b[30]), .Z(n1346) );
  CENX1 U1901 ( .A(n1711), .B(n109), .Z(n1095) );
  CEOX1 U1902 ( .A(n825), .B(n839), .Z(n382) );
  CENX1 U1903 ( .A(n1706), .B(n104), .Z(n1098) );
  CNR2X1 U1904 ( .A(n1615), .B(n1614), .Z(n280) );
  CENX1 U1905 ( .A(n1724), .B(n1391), .Z(n1325) );
  CENX1 U1906 ( .A(n1755), .B(n1392), .Z(n1170) );
  CENX1 U1907 ( .A(n1707), .B(n1400), .Z(n1114) );
  CENX1 U1908 ( .A(n1723), .B(b[29]), .Z(n1314) );
  CENX1 U1909 ( .A(n1702), .B(n109), .Z(n1093) );
  CENX1 U1910 ( .A(n1711), .B(n113), .Z(n1090) );
  CENX1 U1911 ( .A(n1709), .B(n113), .Z(n1091) );
  CENX1 U1912 ( .A(n1740), .B(n1388), .Z(n1235) );
  CENX1 U1913 ( .A(n1748), .B(n1389), .Z(n1211) );
  CENX1 U1914 ( .A(n1748), .B(n1390), .Z(n1212) );
  CENX1 U1915 ( .A(n1740), .B(n1389), .Z(n1236) );
  CENX1 U1916 ( .A(n1740), .B(n1386), .Z(n1233) );
  CENX1 U1917 ( .A(n1748), .B(n1388), .Z(n1210) );
  CENX1 U1918 ( .A(n1709), .B(n104), .Z(n1103) );
  CENX1 U1919 ( .A(n1709), .B(n109), .Z(n1096) );
  CENX1 U1920 ( .A(a[10]), .B(n1749), .Z(n1611) );
  CIVX2 U1921 ( .A(n12), .Z(n1727) );
  CEOXL U1922 ( .A(a[26]), .B(n104), .Z(n1412) );
  CNIVX2 U1923 ( .A(n1408), .Z(n1711) );
  CNIVX1 U1924 ( .A(n1408), .Z(n1712) );
  CIVX2 U1925 ( .A(n1406), .Z(n1701) );
  CIVX2 U1926 ( .A(n1407), .Z(n1699) );
  CNIVX2 U1927 ( .A(n116), .Z(n1710) );
  CNIVX4 U1928 ( .A(n99), .Z(n1708) );
  CEOXL U1929 ( .A(a[28]), .B(n109), .Z(n1411) );
  CIVX2 U1930 ( .A(n1405), .Z(n1703) );
  CIVX2 U1931 ( .A(n1404), .Z(n1705) );
  CND2X1 U1932 ( .A(n1410), .B(n114), .Z(n115) );
  CEOXL U1933 ( .A(a[30]), .B(a[31]), .Z(n1410) );
  CENX1 U1934 ( .A(n1749), .B(n1395), .Z(n1217) );
  COND2X1 U1935 ( .A(n77), .B(n1160), .C(n1159), .D(n74), .Z(n881) );
  CNR2IX1 U1936 ( .B(n1710), .A(n105), .Z(n830) );
  COND2XL U1937 ( .A(n18), .B(n1315), .C(n1314), .D(n15), .Z(n1029) );
  COND2XL U1938 ( .A(n18), .B(n1343), .C(n1342), .D(n15), .Z(n1057) );
  COND2XL U1939 ( .A(n18), .B(n1341), .C(n1340), .D(n15), .Z(n1055) );
  COND2XL U1940 ( .A(n18), .B(n1338), .C(n1337), .D(n15), .Z(n1052) );
  COND2XL U1941 ( .A(n18), .B(n1316), .C(n1315), .D(n15), .Z(n1030) );
  COND2XL U1942 ( .A(n18), .B(n1339), .C(n1338), .D(n15), .Z(n1053) );
  COND2XL U1943 ( .A(n18), .B(n1336), .C(n1335), .D(n15), .Z(n1050) );
  COND2XL U1944 ( .A(n18), .B(n1335), .C(n1334), .D(n15), .Z(n1049) );
  COND2XL U1945 ( .A(n18), .B(n1337), .C(n1336), .D(n15), .Z(n1051) );
  COND2XL U1946 ( .A(n18), .B(n1332), .C(n1331), .D(n15), .Z(n1046) );
  COND2XL U1947 ( .A(n18), .B(n1327), .C(n1326), .D(n15), .Z(n1041) );
  COND2XL U1948 ( .A(n18), .B(n1318), .C(n1317), .D(n15), .Z(n1032) );
  CENX1 U1949 ( .A(n1742), .B(n1396), .Z(n1243) );
  CENX1 U1950 ( .A(n1748), .B(n1396), .Z(n1218) );
  COND2X1 U1951 ( .A(n53), .B(n1220), .C(n1219), .D(n1583), .Z(n938) );
  COND2X1 U1952 ( .A(n53), .B(n1226), .C(n1225), .D(n1583), .Z(n944) );
  COND2X1 U1953 ( .A(n53), .B(n1227), .C(n1226), .D(n1583), .Z(n945) );
  COND2XL U1954 ( .A(n97), .B(n1115), .C(n1114), .D(n95), .Z(n839) );
  COND2XL U1955 ( .A(n97), .B(n1117), .C(n1116), .D(n95), .Z(n841) );
  COND2XL U1956 ( .A(n1123), .B(n97), .C(n95), .D(n1122), .Z(n847) );
  COND2XL U1957 ( .A(n97), .B(n1118), .C(n1117), .D(n95), .Z(n842) );
  CND2IXL U1958 ( .B(n1710), .A(n86), .Z(n1137) );
  CENXL U1959 ( .A(n1735), .B(n1398), .Z(n1272) );
  CENX1 U1960 ( .A(n1761), .B(n1398), .Z(n1157) );
  CFA1XL U1961 ( .A(n850), .B(n952), .CI(n876), .CO(n405), .S(n406) );
  CEO3X1 U1962 ( .A(n1006), .B(n537), .C(n1034), .Z(n506) );
  CND2XL U1963 ( .A(n1006), .B(n537), .Z(n1687) );
  CND2XL U1964 ( .A(n1006), .B(n1034), .Z(n1688) );
  CND2XL U1965 ( .A(n537), .B(n1034), .Z(n1689) );
  CND3XL U1966 ( .A(n1687), .B(n1688), .C(n1689), .Z(n505) );
  CND2XL U1967 ( .A(n484), .B(n486), .Z(n1690) );
  CND2XL U1968 ( .A(n484), .B(n505), .Z(n1691) );
  CND2XL U1969 ( .A(n486), .B(n505), .Z(n1692) );
  CIVX2 U1970 ( .A(n1746), .Z(n1741) );
  COND2XL U1971 ( .A(n44), .B(n1234), .C(n1233), .D(n1582), .Z(n951) );
  COND2XL U1972 ( .A(n1256), .B(n44), .C(n1255), .D(n1582), .Z(n973) );
  CNR2IXL U1973 ( .B(n1710), .A(n1582), .Z(n974) );
  COND2XL U1974 ( .A(n44), .B(n1745), .C(n1582), .D(n1257), .Z(n814) );
  COND2XL U1975 ( .A(n44), .B(n1251), .C(n1250), .D(n1582), .Z(n968) );
  COND2XL U1976 ( .A(n44), .B(n1237), .C(n1236), .D(n1582), .Z(n954) );
  COND2XL U1977 ( .A(n44), .B(n1253), .C(n1252), .D(n1582), .Z(n970) );
  COND2XL U1978 ( .A(n44), .B(n1236), .C(n1235), .D(n1582), .Z(n953) );
  COND2XL U1979 ( .A(n44), .B(n1248), .C(n1247), .D(n1582), .Z(n965) );
  COND2XL U1980 ( .A(n44), .B(n1250), .C(n1249), .D(n1582), .Z(n967) );
  COND2XL U1981 ( .A(n44), .B(n1252), .C(n1251), .D(n1582), .Z(n969) );
  COND2XL U1982 ( .A(n44), .B(n1235), .C(n1234), .D(n1582), .Z(n952) );
  CENX1 U1983 ( .A(n1758), .B(n1394), .Z(n1172) );
  CENX1 U1984 ( .A(n1709), .B(n1758), .Z(n1187) );
  CIVX1 U1985 ( .A(n1759), .Z(n1758) );
  CIVX2 U1986 ( .A(n1762), .Z(n1761) );
  COND2X1 U1987 ( .A(n61), .B(n1199), .C(n1198), .D(n1549), .Z(n918) );
  CENXL U1988 ( .A(n1716), .B(n1398), .Z(n1365) );
  CIVXL U1989 ( .A(n39), .Z(n1745) );
  CENX1 U1990 ( .A(n1740), .B(n1387), .Z(n1234) );
  CEOXL U1991 ( .A(n329), .B(n147), .Z(product[3]) );
  CNR2X1 U1992 ( .A(n248), .B(n251), .Z(n246) );
  COND2XL U1993 ( .A(n18), .B(n1727), .C(n1344), .D(n15), .Z(n817) );
  CENX1 U1994 ( .A(n1725), .B(n1395), .Z(n1329) );
  CFA1XL U1995 ( .A(n854), .B(n956), .CI(n880), .CO(n511), .S(n512) );
  CFA1XL U1996 ( .A(n922), .B(n964), .CI(n1072), .CO(n671), .S(n672) );
  CIVXL U1997 ( .A(n39), .Z(n1747) );
  CIVX1 U1998 ( .A(n1747), .Z(n1742) );
  COND2X1 U1999 ( .A(n77), .B(n1158), .C(n1157), .D(n74), .Z(n879) );
  COND2XL U2000 ( .A(n18), .B(n1320), .C(n1319), .D(n15), .Z(n1034) );
  CND2IXL U2001 ( .B(n1710), .A(n1749), .Z(n1232) );
  CENX1 U2002 ( .A(n1749), .B(n1398), .Z(n1220) );
  CENX1 U2003 ( .A(n1749), .B(n1397), .Z(n1219) );
  CIVX1 U2004 ( .A(n202), .Z(n344) );
  COND2XL U2005 ( .A(n44), .B(n1246), .C(n1245), .D(n1582), .Z(n963) );
  CENXL U2006 ( .A(n1765), .B(n1398), .Z(n1140) );
  CENXL U2007 ( .A(n1765), .B(n1400), .Z(n1142) );
  CIVX1 U2008 ( .A(n1768), .Z(n1766) );
  CFA1XL U2009 ( .A(n908), .B(n946), .CI(n926), .CO(n729), .S(n730) );
  CND3X1 U2010 ( .A(n1696), .B(n1697), .C(n1698), .Z(n583) );
  COND2X1 U2011 ( .A(n69), .B(n1182), .C(n1181), .D(n66), .Z(n902) );
  CENX1 U2012 ( .A(n1740), .B(n1390), .Z(n1237) );
  COND2XL U2013 ( .A(n36), .B(n1738), .C(n33), .D(n1284), .Z(n815) );
  CND2IXL U2014 ( .B(n1710), .A(n1734), .Z(n1284) );
  CIVX1 U2015 ( .A(n1738), .Z(n1734) );
  CND2IXL U2016 ( .B(n1710), .A(n1719), .Z(n1344) );
  COND2XL U2017 ( .A(n18), .B(n1325), .C(n1324), .D(n15), .Z(n1039) );
  COND2XL U2018 ( .A(n61), .B(n1190), .C(n1189), .D(n1549), .Z(n909) );
  COND2XL U2019 ( .A(n61), .B(n1191), .C(n1190), .D(n1550), .Z(n910) );
  CNR2IXL U2020 ( .B(n1710), .A(n1550), .Z(n928) );
  COND2XL U2021 ( .A(n61), .B(n1192), .C(n1191), .D(n1550), .Z(n911) );
  COND2XL U2022 ( .A(n61), .B(n1193), .C(n1192), .D(n1550), .Z(n912) );
  COND2XL U2023 ( .A(n1208), .B(n61), .C(n1207), .D(n1549), .Z(n927) );
  COND2XL U2024 ( .A(n61), .B(n1204), .C(n1203), .D(n1550), .Z(n923) );
  COND2XL U2025 ( .A(n61), .B(n1753), .C(n1550), .D(n1209), .Z(n812) );
  COND2XL U2026 ( .A(n61), .B(n1198), .C(n1197), .D(n1550), .Z(n917) );
  COND2XL U2027 ( .A(n61), .B(n1205), .C(n1204), .D(n1549), .Z(n924) );
  COND2XL U2028 ( .A(n61), .B(n1195), .C(n1194), .D(n1549), .Z(n914) );
  COND2XL U2029 ( .A(n61), .B(n1201), .C(n1200), .D(n1549), .Z(n920) );
  COND2XL U2030 ( .A(n61), .B(n1203), .C(n1202), .D(n1549), .Z(n922) );
  COND2XL U2031 ( .A(n61), .B(n1206), .C(n1205), .D(n1549), .Z(n925) );
  COND2XL U2032 ( .A(n61), .B(n1207), .C(n1206), .D(n1549), .Z(n926) );
  CENX1 U2033 ( .A(n1757), .B(n1393), .Z(n1171) );
  CENX1 U2034 ( .A(n1757), .B(n1395), .Z(n1173) );
  CIVX1 U2035 ( .A(n1759), .Z(n1757) );
  CFA1X1 U2036 ( .A(n853), .B(n955), .CI(n879), .CO(n485), .S(n486) );
  CENXL U2037 ( .A(n1716), .B(n1400), .Z(n1367) );
  CENXL U2038 ( .A(n86), .B(n1400), .Z(n1127) );
  CENX1 U2039 ( .A(n1740), .B(n1400), .Z(n1247) );
  CENXL U2040 ( .A(n1735), .B(n1400), .Z(n1274) );
  CENXL U2041 ( .A(n1751), .B(n1400), .Z(n1199) );
  COND2X1 U2042 ( .A(n77), .B(n1163), .C(n1162), .D(n74), .Z(n884) );
  COND2XL U2043 ( .A(n69), .B(n1759), .C(n66), .D(n1188), .Z(n811) );
  CENXL U2044 ( .A(n1754), .B(n1398), .Z(n1176) );
  CIVX1 U2045 ( .A(n1738), .Z(n1737) );
  COND2X1 U2046 ( .A(n77), .B(n1164), .C(n1163), .D(n74), .Z(n885) );
  CND2IXL U2047 ( .B(n1710), .A(n1728), .Z(n1313) );
  CIVXL U2048 ( .A(n156), .Z(n154) );
  CIVX2 U2049 ( .A(n79), .Z(n1768) );
  CIVXL U2050 ( .A(n1566), .Z(n244) );
  COND1XL U2051 ( .A(n251), .B(n264), .C(n252), .Z(n250) );
  CENX1 U2052 ( .A(n1760), .B(n1400), .Z(n1159) );
  CEOXL U2053 ( .A(n313), .B(n143), .Z(product[7]) );
  CEOXL U2054 ( .A(n321), .B(n145), .Z(product[5]) );
  CEOXL U2055 ( .A(n119), .B(n152), .Z(product[31]) );
  COND2XL U2056 ( .A(n53), .B(n1211), .C(n1210), .D(n1583), .Z(n929) );
  COND2XL U2057 ( .A(n53), .B(n1212), .C(n1211), .D(n1583), .Z(n930) );
  COND2XL U2058 ( .A(n53), .B(n1214), .C(n1213), .D(n1583), .Z(n932) );
  COND2XL U2059 ( .A(n53), .B(n1224), .C(n1223), .D(n1583), .Z(n942) );
  COND2XL U2060 ( .A(n53), .B(n1213), .C(n1212), .D(n1583), .Z(n931) );
  COND2XL U2061 ( .A(n53), .B(n1219), .C(n1218), .D(n1583), .Z(n937) );
  COND2XL U2062 ( .A(n53), .B(n1225), .C(n1224), .D(n1583), .Z(n943) );
  COND2XL U2063 ( .A(n53), .B(n1750), .C(n1583), .D(n1232), .Z(n813) );
  COND2XL U2064 ( .A(n1231), .B(n53), .C(n1230), .D(n1583), .Z(n949) );
  COND2XL U2065 ( .A(n53), .B(n1229), .C(n1228), .D(n1583), .Z(n947) );
  COND2XL U2066 ( .A(n53), .B(n1215), .C(n1214), .D(n1583), .Z(n933) );
  COND2XL U2067 ( .A(n53), .B(n1228), .C(n1227), .D(n1583), .Z(n946) );
  CND2XL U2068 ( .A(n1639), .B(n1637), .Z(n1693) );
  CND2X1 U2069 ( .A(n1639), .B(n1638), .Z(n1694) );
  CND2XL U2070 ( .A(n1637), .B(n1638), .Z(n1695) );
  CND3X1 U2071 ( .A(n1693), .B(n1694), .C(n1695), .Z(n603) );
  CND2XL U2072 ( .A(n340), .B(n172), .Z(n122) );
  CND2XL U2073 ( .A(n1642), .B(n1640), .Z(n1696) );
  CND2X1 U2074 ( .A(n1642), .B(n1641), .Z(n1697) );
  CND2XL U2075 ( .A(n1640), .B(n1641), .Z(n1698) );
  COND2XL U2076 ( .A(n69), .B(n1171), .C(n1170), .D(n66), .Z(n891) );
  COND2XL U2077 ( .A(n69), .B(n1172), .C(n1171), .D(n66), .Z(n892) );
  COND2XL U2078 ( .A(n1187), .B(n69), .C(n1186), .D(n66), .Z(n907) );
  COND2XL U2079 ( .A(n69), .B(n1174), .C(n1173), .D(n66), .Z(n894) );
  COND2XL U2080 ( .A(n69), .B(n1185), .C(n1184), .D(n66), .Z(n905) );
  CND2X1 U2081 ( .A(n440), .B(n465), .Z(n172) );
  COAN1X1 U2082 ( .A(n212), .B(n202), .C(n203), .Z(n199) );
  CNR2X1 U2083 ( .A(n171), .B(n176), .Z(n169) );
  COND2XL U2084 ( .A(n27), .B(n1286), .C(n1285), .D(n24), .Z(n1001) );
  COND2XL U2085 ( .A(n27), .B(n1288), .C(n1287), .D(n24), .Z(n1003) );
  COND2XL U2086 ( .A(n27), .B(n1287), .C(n1286), .D(n24), .Z(n1002) );
  COND2XL U2087 ( .A(n27), .B(n1299), .C(n1298), .D(n24), .Z(n1014) );
  COND2XL U2088 ( .A(n27), .B(n1305), .C(n1304), .D(n24), .Z(n1020) );
  COND2XL U2089 ( .A(n27), .B(n1307), .C(n1306), .D(n24), .Z(n1022) );
  COND2XL U2090 ( .A(n27), .B(n1300), .C(n1299), .D(n24), .Z(n1015) );
  COND2XL U2091 ( .A(n27), .B(n1289), .C(n1288), .D(n24), .Z(n1004) );
  COND2XL U2092 ( .A(n27), .B(n1309), .C(n1308), .D(n24), .Z(n1024) );
  COND2XL U2093 ( .A(n27), .B(n1294), .C(n1293), .D(n24), .Z(n1009) );
  COND2XL U2094 ( .A(n27), .B(n1297), .C(n1296), .D(n24), .Z(n1012) );
  COND2XL U2095 ( .A(n27), .B(n1310), .C(n1309), .D(n24), .Z(n1025) );
  COND2XL U2096 ( .A(n27), .B(n1303), .C(n1302), .D(n24), .Z(n1018) );
  COND2XL U2097 ( .A(n27), .B(n1308), .C(n1307), .D(n24), .Z(n1023) );
  COND2XL U2098 ( .A(n27), .B(n1291), .C(n1290), .D(n24), .Z(n1006) );
  COND2XL U2099 ( .A(n27), .B(n1304), .C(n1303), .D(n24), .Z(n1019) );
  COND2XL U2100 ( .A(n27), .B(n1296), .C(n1295), .D(n24), .Z(n1011) );
  CNR2IXL U2101 ( .B(n1710), .A(n24), .Z(n1028) );
  COND2XL U2102 ( .A(n27), .B(n1293), .C(n1292), .D(n24), .Z(n1008) );
  COND2XL U2103 ( .A(n27), .B(n1295), .C(n1294), .D(n24), .Z(n1010) );
  COND2XL U2104 ( .A(n27), .B(n1301), .C(n1300), .D(n24), .Z(n1016) );
  COND2XL U2105 ( .A(n27), .B(n1302), .C(n1301), .D(n24), .Z(n1017) );
  COND2XL U2106 ( .A(n27), .B(n1298), .C(n1297), .D(n24), .Z(n1013) );
  COND2XL U2107 ( .A(n27), .B(n1312), .C(n1311), .D(n24), .Z(n1027) );
  COND2XL U2108 ( .A(n27), .B(n1733), .C(n24), .D(n1313), .Z(n816) );
  COND2XL U2109 ( .A(n27), .B(n1311), .C(n1310), .D(n24), .Z(n1026) );
  CENXL U2110 ( .A(n1723), .B(n1398), .Z(n1332) );
  COND2XL U2111 ( .A(n77), .B(n1154), .C(n1153), .D(n74), .Z(n875) );
  COND2XL U2112 ( .A(n1168), .B(n77), .C(n1167), .D(n74), .Z(n889) );
  COND2XL U2113 ( .A(n77), .B(n1156), .C(n1155), .D(n74), .Z(n877) );
  COND2XL U2114 ( .A(n77), .B(n1155), .C(n1154), .D(n74), .Z(n876) );
  CNR2IXL U2115 ( .B(n1710), .A(n74), .Z(n890) );
  COND2XL U2116 ( .A(n77), .B(n1166), .C(n1165), .D(n74), .Z(n887) );
  COND2XL U2117 ( .A(n77), .B(n1762), .C(n74), .D(n1169), .Z(n810) );
  COND2XL U2118 ( .A(n77), .B(n1162), .C(n1161), .D(n74), .Z(n883) );
  CND2IXL U2119 ( .B(n1710), .A(n1757), .Z(n1188) );
  COND2XL U2120 ( .A(n77), .B(n1165), .C(n1164), .D(n74), .Z(n886) );
  CND2X4 U2121 ( .A(n1422), .B(n33), .Z(n36) );
  CIVXL U2122 ( .A(n1727), .Z(n1719) );
  CIVXL U2123 ( .A(n1727), .Z(n1720) );
  CIVXL U2124 ( .A(n1727), .Z(n1721) );
  CIVXL U2125 ( .A(n1727), .Z(n1722) );
  CIVXL U2126 ( .A(n1727), .Z(n1724) );
  CIVXL U2127 ( .A(n1727), .Z(n1725) );
  CIVXL U2128 ( .A(n1727), .Z(n1726) );
  CIVXL U2129 ( .A(n1733), .Z(n1728) );
  CIVXL U2130 ( .A(n1733), .Z(n1731) );
  CIVXL U2131 ( .A(n1733), .Z(n1732) );
  CIVXL U2132 ( .A(n1747), .Z(n1743) );
  CIVXL U2133 ( .A(n1747), .Z(n1744) );
  CIVXL U2134 ( .A(n1759), .Z(n1755) );
  CIVXL U2135 ( .A(n1759), .Z(n1756) );
  CIVXL U2136 ( .A(n1768), .Z(n1764) );
  CIVXL U2137 ( .A(n1768), .Z(n1765) );
  CIVX2 U2138 ( .A(n149), .Z(product[1]) );
  CIVX2 U2139 ( .A(n289), .Z(n357) );
  CIVX2 U2140 ( .A(n1682), .Z(n356) );
  CIVX2 U2141 ( .A(n275), .Z(n354) );
  CIVX2 U2142 ( .A(n248), .Z(n350) );
  CIVX2 U2143 ( .A(n187), .Z(n342) );
  CIVX2 U2144 ( .A(n336), .Z(n334) );
  CIVX2 U2145 ( .A(n333), .Z(n331) );
  CIVX2 U2146 ( .A(n325), .Z(n323) );
  CIVX2 U2147 ( .A(n317), .Z(n315) );
  CIVX2 U2148 ( .A(n309), .Z(n307) );
  CIVX2 U2149 ( .A(n1679), .Z(n301) );
  CIVX2 U2150 ( .A(n1680), .Z(n296) );
  CIVX2 U2151 ( .A(n292), .Z(n291) );
  CIVX2 U2152 ( .A(n283), .Z(n282) );
  CIVX2 U2153 ( .A(n281), .Z(n279) );
  CIVX2 U2154 ( .A(n280), .Z(n355) );
  CIVX2 U2155 ( .A(n271), .Z(n269) );
  CIVX2 U2156 ( .A(n259), .Z(n261) );
  CIVX2 U2157 ( .A(n258), .Z(n352) );
  CIVX2 U2158 ( .A(n243), .Z(n241) );
  CIVX2 U2159 ( .A(n238), .Z(n236) );
  CIVX2 U2160 ( .A(n225), .Z(n347) );
  CIVX2 U2161 ( .A(n214), .Z(n216) );
  CIVX2 U2162 ( .A(n212), .Z(n210) );
  CIVX2 U2163 ( .A(n193), .Z(n191) );
  CIVX2 U2164 ( .A(n192), .Z(n343) );
  CIVX2 U2165 ( .A(n182), .Z(n184) );
  CIVX2 U2166 ( .A(n165), .Z(n163) );
  CIVX2 U2167 ( .A(n160), .Z(n158) );
  CIVX2 U2168 ( .A(n86), .Z(n1440) );
  CIVX2 U2169 ( .A(n1708), .Z(n1438) );
  CIVX2 U2170 ( .A(n104), .Z(n1437) );
  CIVX2 U2171 ( .A(n109), .Z(n1436) );
  CIVX2 U2172 ( .A(n113), .Z(n1435) );
endmodule


module calc_DW02_mult_2_stage_6 ( A, B, TC, CLK, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC, CLK;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, \A_extended[32] ,
         \B_extended[32] , n6, n8, n10, n12, n14, n16, n17, n20, n21, n22, n23,
         n24;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33;
  assign \A_extended[32]  = A[31];
  assign \B_extended[32]  = B[31];

  calc_DW_mult_tc_15 mult_96 ( .a({\A_extended[32] , \A_extended[32] , A[30:0]}), .b({\B_extended[32] , \B_extended[32] , B[30:0]}), .product({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, PRODUCT[31:9], n26, 
        n27, n28, n29, n30, n31, n32, n33, n34}), .i_retiming_group_1_clk(CLK)
         );
  CFD1QXL clk_r_REG272_S1 ( .D(n30), .CP(CLK), .Q(n21) );
  CFD1QXL clk_r_REG266_S1 ( .D(n26), .CP(CLK), .Q(PRODUCT[8]) );
  CFD1QXL clk_r_REG268_S1 ( .D(n27), .CP(CLK), .Q(n24) );
  CFD1QXL clk_r_REG270_S1 ( .D(n28), .CP(CLK), .Q(n23) );
  CFD1QXL clk_r_REG271_S1 ( .D(n29), .CP(CLK), .Q(n22) );
  CFD1QXL clk_r_REG273_S1 ( .D(n31), .CP(CLK), .Q(n20) );
  CFD1QXL clk_r_REG276_S1 ( .D(n34), .CP(CLK), .Q(n17) );
  CFD1QXL clk_r_REG274_S1 ( .D(n32), .CP(CLK), .Q(PRODUCT[2]) );
  CFD1QXL clk_r_REG275_S1 ( .D(n33), .CP(CLK), .Q(PRODUCT[1]) );
  CNIVX1 U1 ( .A(n6), .Z(PRODUCT[0]) );
  CNIVX1 U2 ( .A(n17), .Z(n6) );
  CNIVX1 U3 ( .A(n8), .Z(PRODUCT[4]) );
  CNIVX1 U4 ( .A(n21), .Z(n8) );
  CNIVX1 U5 ( .A(n10), .Z(PRODUCT[5]) );
  CNIVX1 U6 ( .A(n22), .Z(n10) );
  CNIVX1 U7 ( .A(n12), .Z(PRODUCT[3]) );
  CNIVX1 U8 ( .A(n20), .Z(n12) );
  CNIVX1 U9 ( .A(n14), .Z(PRODUCT[7]) );
  CNIVX1 U10 ( .A(n24), .Z(n14) );
  CNIVX1 U11 ( .A(n16), .Z(PRODUCT[6]) );
  CNIVX1 U12 ( .A(n23), .Z(n16) );
endmodule


module calc ( clk, rst, A, B, C, pushA, stopA, pushB, stopB, pushC, stopC, Z, 
        pushZ );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  output [31:0] Z;
  input clk, rst, pushA, pushB, pushC;
  output stopA, stopB, stopC, pushZ;
  wire   all_in, all_in1, all_in2, all_in3, all_in4, all_in5, all_in6, all_in7,
         all_in8, all_in9, N7, n13, n14, n15, n16, n18, n20, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, \w9[0] ,
         \w9[10] , \w9[11] , \w9[12] , \w9[13] , \w9[14] , \w9[15] , \w9[16] ,
         \w9[17] , \w9[18] , \w9[19] , \w9[1] , \w9[20] , \w9[21] , \w9[22] ,
         \w9[23] , \w9[24] , \w9[25] , \w9[26] , \w9[27] , \w9[28] , \w9[29] ,
         \w9[2] , \w9[30] , \w9[31] , \w9[3] , \w9[4] , \w9[5] , \w9[6] ,
         \w9[7] , \w9[8] , \w9[9] , \w10[0] , \w10[10] , \w10[11] , \w10[12] ,
         \w10[13] , \w10[14] , \w10[15] , \w10[16] , \w10[17] , \w10[18] ,
         \w10[19] , \w10[1] , \w10[20] , \w10[21] , \w10[22] , \w10[23] ,
         \w10[24] , \w10[25] , \w10[26] , \w10[27] , \w10[28] , \w10[29] ,
         \w10[2] , \w10[30] , \w10[31] , \w10[3] , \w10[4] , \w10[5] ,
         \w10[6] , \w10[7] , \w10[8] , \w10[9] , n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526;
  wire   [63:0] w1;
  wire   [63:0] w2;
  wire   [63:0] w3;
  wire   [63:0] w4;
  wire   [63:0] w5;
  wire   [63:0] w6;
  wire   [63:0] w7;
  wire   [63:0] w8;
  wire   [63:0] w11;
  wire   [31:0] captA;
  wire   [31:0] captB;
  wire   [31:0] captC;
  wire   [31:0] f01;
  wire   [31:0] f02;
  wire   [31:0] f03;
  wire   [31:0] f11;
  wire   [31:0] f12;
  wire   [31:0] f13;
  wire   [31:0] f14;
  wire   [31:0] f15;
  wire   [31:0] f21;
  wire   [31:0] f23;
  wire   [31:0] f26;
  wire   [31:0] f27;
  wire   [31:0] f28;
  wire   [31:0] f31;
  wire   [31:0] f32;
  wire   [31:0] f34;
  wire   [31:0] f35;
  wire   [31:0] f36;
  wire   [31:0] f37;
  wire   [31:0] f41;
  wire   [31:0] f42;
  wire   [31:0] f44;
  wire   [31:0] f46;
  wire   [31:0] f51;
  wire   [31:0] f52;
  wire   [31:0] f53;
  wire   [31:0] f54;
  wire   [31:0] f61;
  wire   [31:0] f62;
  wire   [31:0] f63;
  wire   [31:0] f71;
  wire   [31:0] f72;
  wire   [2:0] seen_d;
  wire   [31:0] f38;
  wire   [31:0] s41;
  wire   [31:0] s42;
  wire   [31:0] s54;
  wire   [31:0] s61;
  wire   [31:0] s72;
  wire   [31:0] res_d;
  wire   [31:0] s81;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154, SYNOPSYS_UNCONNECTED__155, 
        SYNOPSYS_UNCONNECTED__156, SYNOPSYS_UNCONNECTED__157, 
        SYNOPSYS_UNCONNECTED__158, SYNOPSYS_UNCONNECTED__159, 
        SYNOPSYS_UNCONNECTED__160, SYNOPSYS_UNCONNECTED__161, 
        SYNOPSYS_UNCONNECTED__162, SYNOPSYS_UNCONNECTED__163, 
        SYNOPSYS_UNCONNECTED__164, SYNOPSYS_UNCONNECTED__165, 
        SYNOPSYS_UNCONNECTED__166, SYNOPSYS_UNCONNECTED__167, 
        SYNOPSYS_UNCONNECTED__168, SYNOPSYS_UNCONNECTED__169, 
        SYNOPSYS_UNCONNECTED__170, SYNOPSYS_UNCONNECTED__171, 
        SYNOPSYS_UNCONNECTED__172, SYNOPSYS_UNCONNECTED__173, 
        SYNOPSYS_UNCONNECTED__174, SYNOPSYS_UNCONNECTED__175, 
        SYNOPSYS_UNCONNECTED__176, SYNOPSYS_UNCONNECTED__177, 
        SYNOPSYS_UNCONNECTED__178, SYNOPSYS_UNCONNECTED__179, 
        SYNOPSYS_UNCONNECTED__180, SYNOPSYS_UNCONNECTED__181, 
        SYNOPSYS_UNCONNECTED__182, SYNOPSYS_UNCONNECTED__183, 
        SYNOPSYS_UNCONNECTED__184, SYNOPSYS_UNCONNECTED__185, 
        SYNOPSYS_UNCONNECTED__186, SYNOPSYS_UNCONNECTED__187, 
        SYNOPSYS_UNCONNECTED__188, SYNOPSYS_UNCONNECTED__189, 
        SYNOPSYS_UNCONNECTED__190, SYNOPSYS_UNCONNECTED__191, 
        SYNOPSYS_UNCONNECTED__192, SYNOPSYS_UNCONNECTED__193, 
        SYNOPSYS_UNCONNECTED__194, SYNOPSYS_UNCONNECTED__195, 
        SYNOPSYS_UNCONNECTED__196, SYNOPSYS_UNCONNECTED__197, 
        SYNOPSYS_UNCONNECTED__198, SYNOPSYS_UNCONNECTED__199, 
        SYNOPSYS_UNCONNECTED__200, SYNOPSYS_UNCONNECTED__201, 
        SYNOPSYS_UNCONNECTED__202, SYNOPSYS_UNCONNECTED__203, 
        SYNOPSYS_UNCONNECTED__204, SYNOPSYS_UNCONNECTED__205, 
        SYNOPSYS_UNCONNECTED__206, SYNOPSYS_UNCONNECTED__207, 
        SYNOPSYS_UNCONNECTED__208, SYNOPSYS_UNCONNECTED__209, 
        SYNOPSYS_UNCONNECTED__210, SYNOPSYS_UNCONNECTED__211, 
        SYNOPSYS_UNCONNECTED__212, SYNOPSYS_UNCONNECTED__213, 
        SYNOPSYS_UNCONNECTED__214, SYNOPSYS_UNCONNECTED__215, 
        SYNOPSYS_UNCONNECTED__216, SYNOPSYS_UNCONNECTED__217, 
        SYNOPSYS_UNCONNECTED__218, SYNOPSYS_UNCONNECTED__219, 
        SYNOPSYS_UNCONNECTED__220, SYNOPSYS_UNCONNECTED__221, 
        SYNOPSYS_UNCONNECTED__222, SYNOPSYS_UNCONNECTED__223, 
        SYNOPSYS_UNCONNECTED__224, SYNOPSYS_UNCONNECTED__225, 
        SYNOPSYS_UNCONNECTED__226, SYNOPSYS_UNCONNECTED__227, 
        SYNOPSYS_UNCONNECTED__228, SYNOPSYS_UNCONNECTED__229, 
        SYNOPSYS_UNCONNECTED__230, SYNOPSYS_UNCONNECTED__231, 
        SYNOPSYS_UNCONNECTED__232, SYNOPSYS_UNCONNECTED__233, 
        SYNOPSYS_UNCONNECTED__234, SYNOPSYS_UNCONNECTED__235, 
        SYNOPSYS_UNCONNECTED__236, SYNOPSYS_UNCONNECTED__237, 
        SYNOPSYS_UNCONNECTED__238, SYNOPSYS_UNCONNECTED__239, 
        SYNOPSYS_UNCONNECTED__240, SYNOPSYS_UNCONNECTED__241, 
        SYNOPSYS_UNCONNECTED__242, SYNOPSYS_UNCONNECTED__243, 
        SYNOPSYS_UNCONNECTED__244, SYNOPSYS_UNCONNECTED__245, 
        SYNOPSYS_UNCONNECTED__246, SYNOPSYS_UNCONNECTED__247, 
        SYNOPSYS_UNCONNECTED__248, SYNOPSYS_UNCONNECTED__249, 
        SYNOPSYS_UNCONNECTED__250, SYNOPSYS_UNCONNECTED__251, 
        SYNOPSYS_UNCONNECTED__252, SYNOPSYS_UNCONNECTED__253, 
        SYNOPSYS_UNCONNECTED__254, SYNOPSYS_UNCONNECTED__255, 
        SYNOPSYS_UNCONNECTED__256, SYNOPSYS_UNCONNECTED__257, 
        SYNOPSYS_UNCONNECTED__258, SYNOPSYS_UNCONNECTED__259, 
        SYNOPSYS_UNCONNECTED__260, SYNOPSYS_UNCONNECTED__261, 
        SYNOPSYS_UNCONNECTED__262, SYNOPSYS_UNCONNECTED__263, 
        SYNOPSYS_UNCONNECTED__264, SYNOPSYS_UNCONNECTED__265, 
        SYNOPSYS_UNCONNECTED__266, SYNOPSYS_UNCONNECTED__267, 
        SYNOPSYS_UNCONNECTED__268, SYNOPSYS_UNCONNECTED__269, 
        SYNOPSYS_UNCONNECTED__270, SYNOPSYS_UNCONNECTED__271, 
        SYNOPSYS_UNCONNECTED__272, SYNOPSYS_UNCONNECTED__273, 
        SYNOPSYS_UNCONNECTED__274, SYNOPSYS_UNCONNECTED__275, 
        SYNOPSYS_UNCONNECTED__276, SYNOPSYS_UNCONNECTED__277, 
        SYNOPSYS_UNCONNECTED__278, SYNOPSYS_UNCONNECTED__279, 
        SYNOPSYS_UNCONNECTED__280, SYNOPSYS_UNCONNECTED__281, 
        SYNOPSYS_UNCONNECTED__282, SYNOPSYS_UNCONNECTED__283, 
        SYNOPSYS_UNCONNECTED__284, SYNOPSYS_UNCONNECTED__285, 
        SYNOPSYS_UNCONNECTED__286, SYNOPSYS_UNCONNECTED__287, 
        SYNOPSYS_UNCONNECTED__288, SYNOPSYS_UNCONNECTED__289, 
        SYNOPSYS_UNCONNECTED__290, SYNOPSYS_UNCONNECTED__291, 
        SYNOPSYS_UNCONNECTED__292, SYNOPSYS_UNCONNECTED__293, 
        SYNOPSYS_UNCONNECTED__294, SYNOPSYS_UNCONNECTED__295, 
        SYNOPSYS_UNCONNECTED__296, SYNOPSYS_UNCONNECTED__297, 
        SYNOPSYS_UNCONNECTED__298, SYNOPSYS_UNCONNECTED__299, 
        SYNOPSYS_UNCONNECTED__300, SYNOPSYS_UNCONNECTED__301, 
        SYNOPSYS_UNCONNECTED__302, SYNOPSYS_UNCONNECTED__303, 
        SYNOPSYS_UNCONNECTED__304, SYNOPSYS_UNCONNECTED__305, 
        SYNOPSYS_UNCONNECTED__306, SYNOPSYS_UNCONNECTED__307, 
        SYNOPSYS_UNCONNECTED__308, SYNOPSYS_UNCONNECTED__309, 
        SYNOPSYS_UNCONNECTED__310, SYNOPSYS_UNCONNECTED__311, 
        SYNOPSYS_UNCONNECTED__312, SYNOPSYS_UNCONNECTED__313, 
        SYNOPSYS_UNCONNECTED__314, SYNOPSYS_UNCONNECTED__315, 
        SYNOPSYS_UNCONNECTED__316, SYNOPSYS_UNCONNECTED__317, 
        SYNOPSYS_UNCONNECTED__318, SYNOPSYS_UNCONNECTED__319, 
        SYNOPSYS_UNCONNECTED__320, SYNOPSYS_UNCONNECTED__321, 
        SYNOPSYS_UNCONNECTED__322, SYNOPSYS_UNCONNECTED__323, 
        SYNOPSYS_UNCONNECTED__324, SYNOPSYS_UNCONNECTED__325, 
        SYNOPSYS_UNCONNECTED__326, SYNOPSYS_UNCONNECTED__327, 
        SYNOPSYS_UNCONNECTED__328, SYNOPSYS_UNCONNECTED__329, 
        SYNOPSYS_UNCONNECTED__330, SYNOPSYS_UNCONNECTED__331, 
        SYNOPSYS_UNCONNECTED__332, SYNOPSYS_UNCONNECTED__333, 
        SYNOPSYS_UNCONNECTED__334, SYNOPSYS_UNCONNECTED__335, 
        SYNOPSYS_UNCONNECTED__336, SYNOPSYS_UNCONNECTED__337, 
        SYNOPSYS_UNCONNECTED__338, SYNOPSYS_UNCONNECTED__339, 
        SYNOPSYS_UNCONNECTED__340, SYNOPSYS_UNCONNECTED__341, 
        SYNOPSYS_UNCONNECTED__342, SYNOPSYS_UNCONNECTED__343, 
        SYNOPSYS_UNCONNECTED__344, SYNOPSYS_UNCONNECTED__345, 
        SYNOPSYS_UNCONNECTED__346, SYNOPSYS_UNCONNECTED__347, 
        SYNOPSYS_UNCONNECTED__348, SYNOPSYS_UNCONNECTED__349, 
        SYNOPSYS_UNCONNECTED__350, SYNOPSYS_UNCONNECTED__351, 
        SYNOPSYS_UNCONNECTED__352, SYNOPSYS_UNCONNECTED__353, 
        SYNOPSYS_UNCONNECTED__354;

  CFD2QX2 \captA_reg[1]  ( .D(n151), .CP(clk), .CD(n1462), .Q(captA[1]) );
  CFD2QX2 \captB_reg[1]  ( .D(n119), .CP(clk), .CD(n1440), .Q(captB[1]) );
  CFD2QX2 \captC_reg[1]  ( .D(n87), .CP(clk), .CD(n1456), .Q(captC[1]) );
  CFD2QX2 \f01_reg[27]  ( .D(n709), .CP(clk), .CD(n1445), .Q(f01[27]) );
  CFD2QX2 \f01_reg[3]  ( .D(n707), .CP(clk), .CD(n1461), .Q(f01[3]) );
  CFD2QX2 \f02_reg[29]  ( .D(n706), .CP(clk), .CD(n1483), .Q(f02[29]) );
  CFD2QX2 \f02_reg[27]  ( .D(n705), .CP(clk), .CD(n1486), .Q(f02[27]) );
  CFD2QX2 \f02_reg[25]  ( .D(n704), .CP(clk), .CD(n1490), .Q(f02[25]) );
  CFD2QX2 \f02_reg[22]  ( .D(n191), .CP(clk), .CD(n1472), .Q(f02[22]) );
  CFD2QX2 \f02_reg[20]  ( .D(n700), .CP(clk), .CD(n1475), .Q(f02[20]) );
  CFD2QX2 \f02_reg[19]  ( .D(n697), .CP(clk), .CD(n1477), .Q(f02[19]) );
  CFD2QX2 \f02_reg[18]  ( .D(n694), .CP(clk), .CD(n1478), .Q(f02[18]) );
  CFD2QX2 \f02_reg[16]  ( .D(n691), .CP(clk), .CD(n1503), .Q(f02[16]) );
  CFD2QX2 \f02_reg[15]  ( .D(n688), .CP(clk), .CD(n1505), .Q(f02[15]) );
  CFD2QX2 \f02_reg[10]  ( .D(n684), .CP(clk), .CD(n1492), .Q(f02[10]) );
  CFD2QX2 \f03_reg[21]  ( .D(n677), .CP(clk), .CD(n1446), .Q(f03[21]) );
  CFD2QX2 \f03_reg[20]  ( .D(n674), .CP(clk), .CD(n1447), .Q(f03[20]) );
  CFD2QX2 \f03_reg[19]  ( .D(n671), .CP(clk), .CD(n1447), .Q(f03[19]) );
  CFD2QX2 \f03_reg[18]  ( .D(n668), .CP(clk), .CD(n1448), .Q(f03[18]) );
  CFD2QX2 \f03_reg[16]  ( .D(n665), .CP(clk), .CD(n1449), .Q(f03[16]) );
  CFD2QX2 \f03_reg[15]  ( .D(n662), .CP(clk), .CD(n1449), .Q(f03[15]) );
  CFD2QX2 \f03_reg[13]  ( .D(n659), .CP(clk), .CD(n1450), .Q(f03[13]) );
  CFD2QX2 \f03_reg[12]  ( .D(n657), .CP(clk), .CD(n1451), .Q(f03[12]) );
  CFD2QX2 \f12_reg[29]  ( .D(w1[29]), .CP(clk), .CD(n1444), .Q(f12[29]) );
  CFD2QX2 \f12_reg[27]  ( .D(w1[27]), .CP(clk), .CD(n1424), .Q(f12[27]) );
  CFD2QX2 \f12_reg[20]  ( .D(w1[20]), .CP(clk), .CD(n1429), .Q(f12[20]) );
  CFD2QX2 \f12_reg[16]  ( .D(w1[16]), .CP(clk), .CD(n1431), .Q(f12[16]) );
  CFD2QX2 \f12_reg[14]  ( .D(w1[14]), .CP(clk), .CD(n1433), .Q(f12[14]) );
  CFD2QX2 \f12_reg[12]  ( .D(w1[12]), .CP(clk), .CD(n1434), .Q(f12[12]) );
  CFD2QX2 \f12_reg[8]  ( .D(w1[8]), .CP(clk), .CD(n1458), .Q(f12[8]) );
  CFD2QX2 \f12_reg[6]  ( .D(w1[6]), .CP(clk), .CD(n1460), .Q(f12[6]) );
  CFD2QX2 \f12_reg[4]  ( .D(w1[4]), .CP(clk), .CD(n1461), .Q(f12[4]) );
  CFD2QX2 \f12_reg[0]  ( .D(w1[0]), .CP(clk), .CD(n1463), .Q(f12[0]) );
  calc_DW02_mult_2_stage_3 dw8 ( .A({f14[31:2], 1'b0, f14[0]}), .B(f13), .TC(
        1'b1), .CLK(clk), .PRODUCT({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, w8[31:0]}) );
  calc_DW02_mult_2_stage_5 dw6 ( .A(f01), .B(f02), .TC(1'b1), .CLK(clk), 
        .PRODUCT({SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, w6[31:0]}) );
  calc_DW02_mult_2_stage_7 dw4 ( .A(f01), .B(f03), .TC(1'b1), .CLK(clk), 
        .PRODUCT({SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, w4[31:0]}) );
  calc_DW02_mult_2_stage_8 dw3 ( .A(captC), .B({captC[31:1], n188}), .TC(1'b1), 
        .CLK(clk), .PRODUCT({SYNOPSYS_UNCONNECTED__96, 
        SYNOPSYS_UNCONNECTED__97, SYNOPSYS_UNCONNECTED__98, 
        SYNOPSYS_UNCONNECTED__99, SYNOPSYS_UNCONNECTED__100, 
        SYNOPSYS_UNCONNECTED__101, SYNOPSYS_UNCONNECTED__102, 
        SYNOPSYS_UNCONNECTED__103, SYNOPSYS_UNCONNECTED__104, 
        SYNOPSYS_UNCONNECTED__105, SYNOPSYS_UNCONNECTED__106, 
        SYNOPSYS_UNCONNECTED__107, SYNOPSYS_UNCONNECTED__108, 
        SYNOPSYS_UNCONNECTED__109, SYNOPSYS_UNCONNECTED__110, 
        SYNOPSYS_UNCONNECTED__111, SYNOPSYS_UNCONNECTED__112, 
        SYNOPSYS_UNCONNECTED__113, SYNOPSYS_UNCONNECTED__114, 
        SYNOPSYS_UNCONNECTED__115, SYNOPSYS_UNCONNECTED__116, 
        SYNOPSYS_UNCONNECTED__117, SYNOPSYS_UNCONNECTED__118, 
        SYNOPSYS_UNCONNECTED__119, SYNOPSYS_UNCONNECTED__120, 
        SYNOPSYS_UNCONNECTED__121, SYNOPSYS_UNCONNECTED__122, 
        SYNOPSYS_UNCONNECTED__123, SYNOPSYS_UNCONNECTED__124, 
        SYNOPSYS_UNCONNECTED__125, SYNOPSYS_UNCONNECTED__126, 
        SYNOPSYS_UNCONNECTED__127, w3[31:2], SYNOPSYS_UNCONNECTED__128, w3[0]}) );
  calc_DW02_mult_2_stage_9 dw2 ( .A(captB), .B({captB[31:1], n680}), .TC(1'b1), 
        .CLK(clk), .PRODUCT({SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154, SYNOPSYS_UNCONNECTED__155, 
        SYNOPSYS_UNCONNECTED__156, SYNOPSYS_UNCONNECTED__157, 
        SYNOPSYS_UNCONNECTED__158, SYNOPSYS_UNCONNECTED__159, 
        SYNOPSYS_UNCONNECTED__160, w2[31:2], SYNOPSYS_UNCONNECTED__161, w2[0]}) );
  calc_DW02_mult_2_stage_10 dw1 ( .A(captA), .B({captA[31:1], n503}), .TC(1'b1), .CLK(clk), .PRODUCT({SYNOPSYS_UNCONNECTED__162, SYNOPSYS_UNCONNECTED__163, 
        SYNOPSYS_UNCONNECTED__164, SYNOPSYS_UNCONNECTED__165, 
        SYNOPSYS_UNCONNECTED__166, SYNOPSYS_UNCONNECTED__167, 
        SYNOPSYS_UNCONNECTED__168, SYNOPSYS_UNCONNECTED__169, 
        SYNOPSYS_UNCONNECTED__170, SYNOPSYS_UNCONNECTED__171, 
        SYNOPSYS_UNCONNECTED__172, SYNOPSYS_UNCONNECTED__173, 
        SYNOPSYS_UNCONNECTED__174, SYNOPSYS_UNCONNECTED__175, 
        SYNOPSYS_UNCONNECTED__176, SYNOPSYS_UNCONNECTED__177, 
        SYNOPSYS_UNCONNECTED__178, SYNOPSYS_UNCONNECTED__179, 
        SYNOPSYS_UNCONNECTED__180, SYNOPSYS_UNCONNECTED__181, 
        SYNOPSYS_UNCONNECTED__182, SYNOPSYS_UNCONNECTED__183, 
        SYNOPSYS_UNCONNECTED__184, SYNOPSYS_UNCONNECTED__185, 
        SYNOPSYS_UNCONNECTED__186, SYNOPSYS_UNCONNECTED__187, 
        SYNOPSYS_UNCONNECTED__188, SYNOPSYS_UNCONNECTED__189, 
        SYNOPSYS_UNCONNECTED__190, SYNOPSYS_UNCONNECTED__191, 
        SYNOPSYS_UNCONNECTED__192, SYNOPSYS_UNCONNECTED__193, w1[31:2], 
        SYNOPSYS_UNCONNECTED__194, w1[0]}) );
  calc_DW01_add_6 add_314 ( .A(f71), .B(f72), .CI(1'b0), .SUM(s81) );
  calc_DW01_add_7 add_311 ( .A(f62), .B(f63), .CI(1'b0), .SUM(s72) );
  calc_DW01_add_8 add_304 ( .A(f51), .B({n1420, f53[30:0]}), .CI(1'b0), .SUM(
        s61) );
  calc_DW01_add_9 add_301 ( .A(f44), .B({f46[31:2], 1'b0, f46[0]}), .CI(1'b0), 
        .SUM(s54) );
  calc_DW01_add_10 add_291 ( .A(f35), .B({n1419, f32[30:0]}), .CI(1'b0), .SUM(
        s42) );
  calc_DW01_add_11 add_290 ( .A(f34), .B(f38), .CI(1'b0), .SUM(s41) );
  CFD2QXL \f13_reg[17]  ( .D(n246), .CP(clk), .CD(n1512), .Q(f13[17]) );
  CFD2QXL \f13_reg[15]  ( .D(n244), .CP(clk), .CD(n1512), .Q(f13[15]) );
  CFD2QXL \f13_reg[19]  ( .D(n242), .CP(clk), .CD(n1512), .Q(f13[19]) );
  CFD2QXL \f13_reg[9]  ( .D(n239), .CP(clk), .CD(n1512), .Q(f13[9]) );
  CFD2QXL \f13_reg[7]  ( .D(n236), .CP(clk), .CD(n1512), .Q(f13[7]) );
  CFD2QX1 \f12_reg[19]  ( .D(w1[19]), .CP(clk), .CD(n1511), .Q(f12[19]) );
  CFD2QXL \f13_reg[3]  ( .D(n233), .CP(clk), .CD(n1512), .Q(f13[3]) );
  CFD2QXL \f27_reg[17]  ( .D(n1417), .CP(clk), .CD(n1512), .Q(f27[17]) );
  CFD2QXL \f27_reg[16]  ( .D(w5[16]), .CP(clk), .CD(n1512), .Q(f27[16]) );
  CFD2QXL \f13_reg[11]  ( .D(n230), .CP(clk), .CD(n1512), .Q(f13[11]) );
  CFD2QX1 \f12_reg[7]  ( .D(w1[7]), .CP(clk), .CD(n1511), .Q(f12[7]) );
  CFD2QXL \f13_reg[12]  ( .D(n229), .CP(clk), .CD(n1512), .Q(f13[12]) );
  CFD2QX1 \f12_reg[3]  ( .D(w1[3]), .CP(clk), .CD(n1510), .Q(f12[3]) );
  CFD2QXL \f27_reg[0]  ( .D(w5[0]), .CP(clk), .CD(n1512), .Q(f27[0]) );
  CFD2QXL \f13_reg[1]  ( .D(n460), .CP(clk), .CD(n1512), .Q(f13[1]) );
  CFD2QX1 \f02_reg[11]  ( .D(n463), .CP(clk), .CD(n1511), .Q(f02[11]) );
  CFD2QX4 \f02_reg[14]  ( .D(n464), .CP(clk), .CD(n1424), .Q(f02[14]) );
  CFD2QXL \f27_reg[2]  ( .D(w5[2]), .CP(clk), .CD(n1512), .Q(f27[2]) );
  CFD2QXL \f27_reg[1]  ( .D(w5[1]), .CP(clk), .CD(n1512), .Q(f27[1]) );
  CFD2QX1 \f12_reg[11]  ( .D(w1[11]), .CP(clk), .CD(n1511), .Q(f12[11]) );
  CFD2QX1 \f12_reg[13]  ( .D(w1[13]), .CP(clk), .CD(n1511), .Q(f12[13]) );
  CFD2QXL \f13_reg[21]  ( .D(n186), .CP(clk), .CD(n1511), .Q(f13[21]) );
  CFD2QX1 \f12_reg[15]  ( .D(w1[15]), .CP(clk), .CD(n1511), .Q(f12[15]) );
  CFD2QX1 \f12_reg[17]  ( .D(w1[17]), .CP(clk), .CD(n1511), .Q(f12[17]) );
  CFD2QXL \f27_reg[4]  ( .D(w5[4]), .CP(clk), .CD(n1512), .Q(f27[4]) );
  CFD2QX1 \f12_reg[21]  ( .D(w1[21]), .CP(clk), .CD(n1510), .Q(f12[21]) );
  CFD2QX1 \f12_reg[9]  ( .D(w1[9]), .CP(clk), .CD(n1511), .Q(f12[9]) );
  CFD2QXL \f13_reg[23]  ( .D(n476), .CP(clk), .CD(n1512), .Q(f13[23]) );
  CFD2QX4 \f03_reg[14]  ( .D(n319), .CP(clk), .CD(n1424), .Q(f03[14]) );
  calc_DW02_mult_2_stage_0 dw11 ( .A({\w10[31] , \w10[30] , \w10[29] , 
        \w10[28] , \w10[27] , \w10[26] , \w10[25] , \w10[24] , \w10[23] , 
        \w10[22] , \w10[21] , \w10[20] , \w10[19] , \w10[18] , \w10[17] , 
        \w10[16] , \w10[15] , \w10[14] , \w10[13] , \w10[12] , \w10[11] , 
        \w10[10] , \w10[9] , \w10[8] , \w10[7] , \w10[6] , \w10[5] , \w10[4] , 
        \w10[3] , \w10[2] , \w10[1] , \w10[0] }), .B(f36), .TC(1'b1), .CLK(clk), .PRODUCT({SYNOPSYS_UNCONNECTED__195, SYNOPSYS_UNCONNECTED__196, 
        SYNOPSYS_UNCONNECTED__197, SYNOPSYS_UNCONNECTED__198, 
        SYNOPSYS_UNCONNECTED__199, SYNOPSYS_UNCONNECTED__200, 
        SYNOPSYS_UNCONNECTED__201, SYNOPSYS_UNCONNECTED__202, 
        SYNOPSYS_UNCONNECTED__203, SYNOPSYS_UNCONNECTED__204, 
        SYNOPSYS_UNCONNECTED__205, SYNOPSYS_UNCONNECTED__206, 
        SYNOPSYS_UNCONNECTED__207, SYNOPSYS_UNCONNECTED__208, 
        SYNOPSYS_UNCONNECTED__209, SYNOPSYS_UNCONNECTED__210, 
        SYNOPSYS_UNCONNECTED__211, SYNOPSYS_UNCONNECTED__212, 
        SYNOPSYS_UNCONNECTED__213, SYNOPSYS_UNCONNECTED__214, 
        SYNOPSYS_UNCONNECTED__215, SYNOPSYS_UNCONNECTED__216, 
        SYNOPSYS_UNCONNECTED__217, SYNOPSYS_UNCONNECTED__218, 
        SYNOPSYS_UNCONNECTED__219, SYNOPSYS_UNCONNECTED__220, 
        SYNOPSYS_UNCONNECTED__221, SYNOPSYS_UNCONNECTED__222, 
        SYNOPSYS_UNCONNECTED__223, SYNOPSYS_UNCONNECTED__224, 
        SYNOPSYS_UNCONNECTED__225, SYNOPSYS_UNCONNECTED__226, w11[31:0]}) );
  calc_DW02_mult_2_stage_1 dw10 ( .A({\w9[31] , \w9[30] , \w9[29] , \w9[28] , 
        \w9[27] , \w9[26] , \w9[25] , \w9[24] , \w9[23] , \w9[22] , \w9[21] , 
        \w9[20] , \w9[19] , \w9[18] , \w9[17] , \w9[16] , \w9[15] , \w9[14] , 
        \w9[13] , \w9[12] , \w9[11] , \w9[10] , \w9[9] , \w9[8] , \w9[7] , 
        \w9[6] , \w9[5] , \w9[4] , \w9[3] , \w9[2] , \w9[1] , \w9[0] }), .B(
        f21), .TC(1'b1), .CLK(clk), .PRODUCT({SYNOPSYS_UNCONNECTED__227, 
        SYNOPSYS_UNCONNECTED__228, SYNOPSYS_UNCONNECTED__229, 
        SYNOPSYS_UNCONNECTED__230, SYNOPSYS_UNCONNECTED__231, 
        SYNOPSYS_UNCONNECTED__232, SYNOPSYS_UNCONNECTED__233, 
        SYNOPSYS_UNCONNECTED__234, SYNOPSYS_UNCONNECTED__235, 
        SYNOPSYS_UNCONNECTED__236, SYNOPSYS_UNCONNECTED__237, 
        SYNOPSYS_UNCONNECTED__238, SYNOPSYS_UNCONNECTED__239, 
        SYNOPSYS_UNCONNECTED__240, SYNOPSYS_UNCONNECTED__241, 
        SYNOPSYS_UNCONNECTED__242, SYNOPSYS_UNCONNECTED__243, 
        SYNOPSYS_UNCONNECTED__244, SYNOPSYS_UNCONNECTED__245, 
        SYNOPSYS_UNCONNECTED__246, SYNOPSYS_UNCONNECTED__247, 
        SYNOPSYS_UNCONNECTED__248, SYNOPSYS_UNCONNECTED__249, 
        SYNOPSYS_UNCONNECTED__250, SYNOPSYS_UNCONNECTED__251, 
        SYNOPSYS_UNCONNECTED__252, SYNOPSYS_UNCONNECTED__253, 
        SYNOPSYS_UNCONNECTED__254, SYNOPSYS_UNCONNECTED__255, 
        SYNOPSYS_UNCONNECTED__256, SYNOPSYS_UNCONNECTED__257, 
        SYNOPSYS_UNCONNECTED__258, \w10[31] , \w10[30] , \w10[29] , \w10[28] , 
        \w10[27] , \w10[26] , \w10[25] , \w10[24] , \w10[23] , \w10[22] , 
        \w10[21] , \w10[20] , \w10[19] , \w10[18] , \w10[17] , \w10[16] , 
        \w10[15] , \w10[14] , \w10[13] , \w10[12] , \w10[11] , \w10[10] , 
        \w10[9] , \w10[8] , \w10[7] , \w10[6] , \w10[5] , \w10[4] , \w10[3] , 
        \w10[2] , \w10[1] , \w10[0] }) );
  calc_DW02_mult_2_stage_2 dw9 ( .A({f12[31:2], 1'b0, f12[0]}), .B(f11), .TC(
        1'b1), .CLK(clk), .PRODUCT({SYNOPSYS_UNCONNECTED__259, 
        SYNOPSYS_UNCONNECTED__260, SYNOPSYS_UNCONNECTED__261, 
        SYNOPSYS_UNCONNECTED__262, SYNOPSYS_UNCONNECTED__263, 
        SYNOPSYS_UNCONNECTED__264, SYNOPSYS_UNCONNECTED__265, 
        SYNOPSYS_UNCONNECTED__266, SYNOPSYS_UNCONNECTED__267, 
        SYNOPSYS_UNCONNECTED__268, SYNOPSYS_UNCONNECTED__269, 
        SYNOPSYS_UNCONNECTED__270, SYNOPSYS_UNCONNECTED__271, 
        SYNOPSYS_UNCONNECTED__272, SYNOPSYS_UNCONNECTED__273, 
        SYNOPSYS_UNCONNECTED__274, SYNOPSYS_UNCONNECTED__275, 
        SYNOPSYS_UNCONNECTED__276, SYNOPSYS_UNCONNECTED__277, 
        SYNOPSYS_UNCONNECTED__278, SYNOPSYS_UNCONNECTED__279, 
        SYNOPSYS_UNCONNECTED__280, SYNOPSYS_UNCONNECTED__281, 
        SYNOPSYS_UNCONNECTED__282, SYNOPSYS_UNCONNECTED__283, 
        SYNOPSYS_UNCONNECTED__284, SYNOPSYS_UNCONNECTED__285, 
        SYNOPSYS_UNCONNECTED__286, SYNOPSYS_UNCONNECTED__287, 
        SYNOPSYS_UNCONNECTED__288, SYNOPSYS_UNCONNECTED__289, 
        SYNOPSYS_UNCONNECTED__290, \w9[31] , \w9[30] , \w9[29] , \w9[28] , 
        \w9[27] , \w9[26] , \w9[25] , \w9[24] , \w9[23] , \w9[22] , \w9[21] , 
        \w9[20] , \w9[19] , \w9[18] , \w9[17] , \w9[16] , \w9[15] , \w9[14] , 
        \w9[13] , \w9[12] , \w9[11] , \w9[10] , \w9[9] , \w9[8] , \w9[7] , 
        \w9[6] , \w9[5] , \w9[4] , \w9[3] , \w9[2] , \w9[1] , \w9[0] }) );
  calc_DW02_mult_2_stage_4 dw7 ( .A({f12[31:10], n1515, f12[8:4], n1518, n1520, 
        1'b0, f12[0]}), .B({w5[31:25], n1421, w5[23], n1423, w5[21:18], n1417, 
        w5[16:0]}), .TC(1'b1), .CLK(clk), .PRODUCT({SYNOPSYS_UNCONNECTED__291, 
        SYNOPSYS_UNCONNECTED__292, SYNOPSYS_UNCONNECTED__293, 
        SYNOPSYS_UNCONNECTED__294, SYNOPSYS_UNCONNECTED__295, 
        SYNOPSYS_UNCONNECTED__296, SYNOPSYS_UNCONNECTED__297, 
        SYNOPSYS_UNCONNECTED__298, SYNOPSYS_UNCONNECTED__299, 
        SYNOPSYS_UNCONNECTED__300, SYNOPSYS_UNCONNECTED__301, 
        SYNOPSYS_UNCONNECTED__302, SYNOPSYS_UNCONNECTED__303, 
        SYNOPSYS_UNCONNECTED__304, SYNOPSYS_UNCONNECTED__305, 
        SYNOPSYS_UNCONNECTED__306, SYNOPSYS_UNCONNECTED__307, 
        SYNOPSYS_UNCONNECTED__308, SYNOPSYS_UNCONNECTED__309, 
        SYNOPSYS_UNCONNECTED__310, SYNOPSYS_UNCONNECTED__311, 
        SYNOPSYS_UNCONNECTED__312, SYNOPSYS_UNCONNECTED__313, 
        SYNOPSYS_UNCONNECTED__314, SYNOPSYS_UNCONNECTED__315, 
        SYNOPSYS_UNCONNECTED__316, SYNOPSYS_UNCONNECTED__317, 
        SYNOPSYS_UNCONNECTED__318, SYNOPSYS_UNCONNECTED__319, 
        SYNOPSYS_UNCONNECTED__320, SYNOPSYS_UNCONNECTED__321, 
        SYNOPSYS_UNCONNECTED__322, w7[31:0]}) );
  calc_DW02_mult_2_stage_6 dw5 ( .A(f02), .B(f03), .TC(1'b1), .CLK(clk), 
        .PRODUCT({SYNOPSYS_UNCONNECTED__323, SYNOPSYS_UNCONNECTED__324, 
        SYNOPSYS_UNCONNECTED__325, SYNOPSYS_UNCONNECTED__326, 
        SYNOPSYS_UNCONNECTED__327, SYNOPSYS_UNCONNECTED__328, 
        SYNOPSYS_UNCONNECTED__329, SYNOPSYS_UNCONNECTED__330, 
        SYNOPSYS_UNCONNECTED__331, SYNOPSYS_UNCONNECTED__332, 
        SYNOPSYS_UNCONNECTED__333, SYNOPSYS_UNCONNECTED__334, 
        SYNOPSYS_UNCONNECTED__335, SYNOPSYS_UNCONNECTED__336, 
        SYNOPSYS_UNCONNECTED__337, SYNOPSYS_UNCONNECTED__338, 
        SYNOPSYS_UNCONNECTED__339, SYNOPSYS_UNCONNECTED__340, 
        SYNOPSYS_UNCONNECTED__341, SYNOPSYS_UNCONNECTED__342, 
        SYNOPSYS_UNCONNECTED__343, SYNOPSYS_UNCONNECTED__344, 
        SYNOPSYS_UNCONNECTED__345, SYNOPSYS_UNCONNECTED__346, 
        SYNOPSYS_UNCONNECTED__347, SYNOPSYS_UNCONNECTED__348, 
        SYNOPSYS_UNCONNECTED__349, SYNOPSYS_UNCONNECTED__350, 
        SYNOPSYS_UNCONNECTED__351, SYNOPSYS_UNCONNECTED__352, 
        SYNOPSYS_UNCONNECTED__353, SYNOPSYS_UNCONNECTED__354, w5[31:0]}) );
  CFD1QXL \res_d_reg[0]  ( .D(n53), .CP(clk), .Q(res_d[0]) );
  CFD1QXL \res_d_reg[1]  ( .D(n52), .CP(clk), .Q(res_d[1]) );
  CFD1QXL \res_d_reg[2]  ( .D(n51), .CP(clk), .Q(res_d[2]) );
  CFD1QXL \res_d_reg[3]  ( .D(n50), .CP(clk), .Q(res_d[3]) );
  CFD1QXL \res_d_reg[4]  ( .D(n49), .CP(clk), .Q(res_d[4]) );
  CFD1QXL \res_d_reg[5]  ( .D(n48), .CP(clk), .Q(res_d[5]) );
  CFD1QXL \res_d_reg[6]  ( .D(n47), .CP(clk), .Q(res_d[6]) );
  CFD1QXL \res_d_reg[7]  ( .D(n46), .CP(clk), .Q(res_d[7]) );
  CFD1QXL \res_d_reg[8]  ( .D(n45), .CP(clk), .Q(res_d[8]) );
  CFD1QXL \res_d_reg[9]  ( .D(n44), .CP(clk), .Q(res_d[9]) );
  CFD1QXL \res_d_reg[10]  ( .D(n43), .CP(clk), .Q(res_d[10]) );
  CFD1QXL \res_d_reg[11]  ( .D(n42), .CP(clk), .Q(res_d[11]) );
  CFD1QXL \res_d_reg[12]  ( .D(n41), .CP(clk), .Q(res_d[12]) );
  CFD1QXL \res_d_reg[13]  ( .D(n40), .CP(clk), .Q(res_d[13]) );
  CFD1QXL \res_d_reg[14]  ( .D(n39), .CP(clk), .Q(res_d[14]) );
  CFD1QXL \res_d_reg[15]  ( .D(n38), .CP(clk), .Q(res_d[15]) );
  CFD1QXL \res_d_reg[16]  ( .D(n37), .CP(clk), .Q(res_d[16]) );
  CFD1QXL \res_d_reg[17]  ( .D(n36), .CP(clk), .Q(res_d[17]) );
  CFD1QXL \res_d_reg[18]  ( .D(n35), .CP(clk), .Q(res_d[18]) );
  CFD1QXL \res_d_reg[19]  ( .D(n34), .CP(clk), .Q(res_d[19]) );
  CFD1QXL \res_d_reg[20]  ( .D(n33), .CP(clk), .Q(res_d[20]) );
  CFD1QXL \res_d_reg[21]  ( .D(n32), .CP(clk), .Q(res_d[21]) );
  CFD1QXL \res_d_reg[22]  ( .D(n31), .CP(clk), .Q(res_d[22]) );
  CFD1QXL \res_d_reg[23]  ( .D(n30), .CP(clk), .Q(res_d[23]) );
  CFD1QXL \res_d_reg[24]  ( .D(n29), .CP(clk), .Q(res_d[24]) );
  CFD1QXL \res_d_reg[25]  ( .D(n28), .CP(clk), .Q(res_d[25]) );
  CFD1QXL \res_d_reg[26]  ( .D(n27), .CP(clk), .Q(res_d[26]) );
  CFD1QXL \res_d_reg[27]  ( .D(n26), .CP(clk), .Q(res_d[27]) );
  CFD1QXL \res_d_reg[28]  ( .D(n25), .CP(clk), .Q(res_d[28]) );
  CFD1QXL \res_d_reg[29]  ( .D(n24), .CP(clk), .Q(res_d[29]) );
  CFD1QXL \res_d_reg[30]  ( .D(n23), .CP(clk), .Q(res_d[30]) );
  CFD1QXL \res_d_reg[31]  ( .D(n22), .CP(clk), .Q(res_d[31]) );
  CFD1QXL \f38_reg[30]  ( .D(n84), .CP(clk), .Q(f38[30]) );
  CFD1QXL \f38_reg[31]  ( .D(n85), .CP(clk), .Q(f38[31]) );
  CFD2QXL \f36_reg[31]  ( .D(n1382), .CP(clk), .CD(n1442), .Q(f36[31]) );
  CFD2QXL \f27_reg[31]  ( .D(w5[31]), .CP(clk), .CD(n1479), .Q(f27[31]) );
  CFD2QXL \f27_reg[30]  ( .D(w5[30]), .CP(clk), .CD(n1481), .Q(f27[30]) );
  CFD2QXL \f27_reg[29]  ( .D(w5[29]), .CP(clk), .CD(n1483), .Q(f27[29]) );
  CFD2QXL \f27_reg[28]  ( .D(w5[28]), .CP(clk), .CD(n1484), .Q(f27[28]) );
  CFD2QXL \f27_reg[27]  ( .D(w5[27]), .CP(clk), .CD(n1486), .Q(f27[27]) );
  CFD2QXL \f27_reg[26]  ( .D(w5[26]), .CP(clk), .CD(n1488), .Q(f27[26]) );
  CFD2QXL \f27_reg[25]  ( .D(w5[25]), .CP(clk), .CD(n1489), .Q(f27[25]) );
  CFD2QXL \f27_reg[24]  ( .D(n1421), .CP(clk), .CD(n1469), .Q(f27[24]) );
  CFD2QXL \f27_reg[23]  ( .D(w5[23]), .CP(clk), .CD(n1470), .Q(f27[23]) );
  CFD2QXL \f27_reg[22]  ( .D(n1423), .CP(clk), .CD(n1472), .Q(f27[22]) );
  CFD2QXL \f27_reg[21]  ( .D(w5[21]), .CP(clk), .CD(n1473), .Q(f27[21]) );
  CFD2QXL \f27_reg[20]  ( .D(w5[20]), .CP(clk), .CD(n1475), .Q(f27[20]) );
  CFD2QXL \f27_reg[19]  ( .D(w5[19]), .CP(clk), .CD(n1476), .Q(f27[19]) );
  CFD2QXL \f27_reg[18]  ( .D(w5[18]), .CP(clk), .CD(n1478), .Q(f27[18]) );
  CFD2QXL \f27_reg[15]  ( .D(w5[15]), .CP(clk), .CD(n1505), .Q(f27[15]) );
  CFD2QXL \f27_reg[14]  ( .D(w5[14]), .CP(clk), .CD(n1506), .Q(f27[14]) );
  CFD2QXL \f27_reg[13]  ( .D(w5[13]), .CP(clk), .CD(n1508), .Q(f27[13]) );
  CFD2QXL \f27_reg[12]  ( .D(w5[12]), .CP(clk), .CD(n1509), .Q(f27[12]) );
  CFD2QXL \f27_reg[11]  ( .D(w5[11]), .CP(clk), .CD(n1490), .Q(f27[11]) );
  CFD2QXL \f27_reg[10]  ( .D(w5[10]), .CP(clk), .CD(n1492), .Q(f27[10]) );
  CFD2QXL \f27_reg[9]  ( .D(w5[9]), .CP(clk), .CD(n1493), .Q(f27[9]) );
  CFD2QXL \f27_reg[8]  ( .D(n1381), .CP(clk), .CD(n1495), .Q(f27[8]) );
  CFD2QXL \f27_reg[7]  ( .D(w5[7]), .CP(clk), .CD(n1497), .Q(f27[7]) );
  CFD2QXL \f27_reg[6]  ( .D(w5[6]), .CP(clk), .CD(n1498), .Q(f27[6]) );
  CFD2QXL \f27_reg[5]  ( .D(w5[5]), .CP(clk), .CD(n1500), .Q(f27[5]) );
  CFD2QXL \f27_reg[3]  ( .D(w5[3]), .CP(clk), .CD(n1436), .Q(f27[3]) );
  CFD2QXL \captA_reg[31]  ( .D(n181), .CP(clk), .CD(n1442), .Q(captA[31]) );
  CFD2QXL \captB_reg[31]  ( .D(n149), .CP(clk), .CD(n1480), .Q(captB[31]) );
  CFD2QXL \captC_reg[31]  ( .D(n117), .CP(clk), .CD(n1464), .Q(captC[31]) );
  CFD1QXL \f38_reg[29]  ( .D(n83), .CP(clk), .Q(f38[29]) );
  CFD1QXL \f38_reg[28]  ( .D(n82), .CP(clk), .Q(f38[28]) );
  CFD2QXL \f34_reg[30]  ( .D(n1368), .CP(clk), .CD(n1443), .Q(f34[30]) );
  CFD2QXL \f35_reg[30]  ( .D(n1370), .CP(clk), .CD(n1481), .Q(f35[30]) );
  CFD2QXL \f44_reg[30]  ( .D(n1372), .CP(clk), .CD(n1481), .Q(f44[30]) );
  CFD2QXL \f51_reg[30]  ( .D(n1374), .CP(clk), .CD(n1481), .Q(f51[30]) );
  CFD2QXL \f62_reg[30]  ( .D(n1376), .CP(clk), .CD(n1480), .Q(f62[30]) );
  CFD2QXL \f46_reg[30]  ( .D(n1364), .CP(clk), .CD(n1465), .Q(f46[30]) );
  CFD2QXL \f53_reg[30]  ( .D(w11[30]), .CP(clk), .CD(n1442), .Q(f53[30]) );
  CFD2QXL \f63_reg[30]  ( .D(n1366), .CP(clk), .CD(n1481), .Q(f63[30]) );
  CFD2QXL \f13_reg[31]  ( .D(f02[31]), .CP(clk), .CD(n1479), .Q(f13[31]) );
  CFD2QXL \f36_reg[30]  ( .D(n1354), .CP(clk), .CD(n1442), .Q(f36[30]) );
  CFD2QXL \f34_reg[31]  ( .D(n1356), .CP(clk), .CD(n1442), .Q(f34[31]) );
  CFD2QXL \f35_reg[31]  ( .D(n1358), .CP(clk), .CD(n1479), .Q(f35[31]) );
  CFD2QXL \f44_reg[31]  ( .D(n1360), .CP(clk), .CD(n1480), .Q(f44[31]) );
  CFD2QXL \f51_reg[31]  ( .D(n1362), .CP(clk), .CD(n1479), .Q(f51[31]) );
  CFD2QXL \f62_reg[31]  ( .D(n1344), .CP(clk), .CD(n1484), .Q(f62[31]) );
  CFD2QXL \f71_reg[31]  ( .D(n1346), .CP(clk), .CD(n1479), .Q(f71[31]) );
  CFD2QXL \f34_reg[29]  ( .D(n1348), .CP(clk), .CD(n1443), .Q(f34[29]) );
  CFD2QXL \f35_reg[29]  ( .D(n1350), .CP(clk), .CD(n1482), .Q(f35[29]) );
  CFD2QXL \f44_reg[29]  ( .D(n1352), .CP(clk), .CD(n1483), .Q(f44[29]) );
  CFD2QXL \f51_reg[29]  ( .D(n1336), .CP(clk), .CD(n1482), .Q(f51[29]) );
  CFD2QXL \f62_reg[29]  ( .D(n1338), .CP(clk), .CD(n1482), .Q(f62[29]) );
  CFD2QXL \f71_reg[30]  ( .D(n1340), .CP(clk), .CD(n1481), .Q(f71[30]) );
  CFD2QXL \f71_reg[29]  ( .D(n1342), .CP(clk), .CD(n1482), .Q(f71[29]) );
  CFD2QXL \f46_reg[31]  ( .D(n1332), .CP(clk), .CD(n1464), .Q(f46[31]) );
  CFD2QXL \f63_reg[31]  ( .D(n1334), .CP(clk), .CD(n1480), .Q(f63[31]) );
  CFD2QXL \f72_reg[31]  ( .D(s72[31]), .CP(clk), .CD(n1490), .Q(f72[31]) );
  CFD2QXL \f32_reg[29]  ( .D(w8[29]), .CP(clk), .CD(n1482), .Q(f32[29]) );
  CFD2QXL \f46_reg[29]  ( .D(n1328), .CP(clk), .CD(n1465), .Q(f46[29]) );
  CFD2QXL \f53_reg[29]  ( .D(w11[29]), .CP(clk), .CD(n1443), .Q(f53[29]) );
  CFD2QXL \f63_reg[29]  ( .D(n1330), .CP(clk), .CD(n1483), .Q(f63[29]) );
  CFD2QXL \f72_reg[30]  ( .D(s72[30]), .CP(clk), .CD(n1480), .Q(f72[30]) );
  CFD2QXL \f72_reg[29]  ( .D(s72[29]), .CP(clk), .CD(n1482), .Q(f72[29]) );
  CFD2QXL \f36_reg[29]  ( .D(n1327), .CP(clk), .CD(n1443), .Q(f36[29]) );
  CFD1QXL \f38_reg[27]  ( .D(n81), .CP(clk), .Q(f38[27]) );
  CFD1QXL \f38_reg[26]  ( .D(n80), .CP(clk), .Q(f38[26]) );
  CFD1QXL \f38_reg[25]  ( .D(n79), .CP(clk), .Q(f38[25]) );
  CFD1QXL \f38_reg[24]  ( .D(n78), .CP(clk), .Q(f38[24]) );
  CFD1QXL \f38_reg[1]  ( .D(n55), .CP(clk), .Q(f38[1]) );
  CFD1QXL \f38_reg[0]  ( .D(n54), .CP(clk), .Q(f38[0]) );
  CFD1QXL \f38_reg[23]  ( .D(n77), .CP(clk), .Q(f38[23]) );
  CFD1QXL \f38_reg[21]  ( .D(n75), .CP(clk), .Q(f38[21]) );
  CFD1QXL \f38_reg[19]  ( .D(n73), .CP(clk), .Q(f38[19]) );
  CFD1QXL \f38_reg[17]  ( .D(n71), .CP(clk), .Q(f38[17]) );
  CFD1QXL \f38_reg[16]  ( .D(n70), .CP(clk), .Q(f38[16]) );
  CFD1QXL \f38_reg[15]  ( .D(n69), .CP(clk), .Q(f38[15]) );
  CFD1QXL \f38_reg[14]  ( .D(n68), .CP(clk), .Q(f38[14]) );
  CFD1QXL \f38_reg[13]  ( .D(n67), .CP(clk), .Q(f38[13]) );
  CFD1QXL \f38_reg[12]  ( .D(n66), .CP(clk), .Q(f38[12]) );
  CFD1QXL \f38_reg[8]  ( .D(n62), .CP(clk), .Q(f38[8]) );
  CFD1QXL \f38_reg[7]  ( .D(n61), .CP(clk), .Q(f38[7]) );
  CFD1QXL \f38_reg[5]  ( .D(n59), .CP(clk), .Q(f38[5]) );
  CFD1QXL \f38_reg[4]  ( .D(n58), .CP(clk), .Q(f38[4]) );
  CFD1QXL \f38_reg[3]  ( .D(n57), .CP(clk), .Q(f38[3]) );
  CFD1QXL \f38_reg[11]  ( .D(n65), .CP(clk), .Q(f38[11]) );
  CFD1QXL \f38_reg[9]  ( .D(n63), .CP(clk), .Q(f38[9]) );
  CFD1QXL \f38_reg[10]  ( .D(n64), .CP(clk), .Q(f38[10]) );
  CFD1QXL \f38_reg[22]  ( .D(n76), .CP(clk), .Q(f38[22]) );
  CFD1QXL \f38_reg[20]  ( .D(n74), .CP(clk), .Q(f38[20]) );
  CFD1QXL \f38_reg[18]  ( .D(n72), .CP(clk), .Q(f38[18]) );
  CFD1QXL \f38_reg[6]  ( .D(n60), .CP(clk), .Q(f38[6]) );
  CFD1QXL \f38_reg[2]  ( .D(n56), .CP(clk), .Q(f38[2]) );
  CFD2QXL \f11_reg[31]  ( .D(f01[31]), .CP(clk), .CD(n1442), .Q(f11[31]) );
  CFD2QXL \f11_reg[30]  ( .D(n1322), .CP(clk), .CD(n1443), .Q(f11[30]) );
  CFD2QXL \f21_reg[31]  ( .D(n1323), .CP(clk), .CD(n1442), .Q(f21[31]) );
  CFD2QXL \f21_reg[30]  ( .D(n1325), .CP(clk), .CD(n1443), .Q(f21[30]) );
  CFD2QXL \f44_reg[1]  ( .D(n1320), .CP(clk), .CD(n1440), .Q(f44[1]) );
  CFD2QXL \f11_reg[29]  ( .D(n1318), .CP(clk), .CD(n1443), .Q(f11[29]) );
  CFD2QXL \f11_reg[28]  ( .D(n1319), .CP(clk), .CD(n1444), .Q(f11[28]) );
  CFD2QXL \f01_reg[25]  ( .D(n1316), .CP(clk), .CD(n1425), .Q(f01[25]) );
  CFD2QXL \captA_reg[30]  ( .D(n180), .CP(clk), .CD(n1443), .Q(captA[30]) );
  CFD2QXL \captA_reg[28]  ( .D(n178), .CP(clk), .CD(n1444), .Q(captA[28]) );
  CFD2QXL \captB_reg[30]  ( .D(n148), .CP(clk), .CD(n1482), .Q(captB[30]) );
  CFD2QXL \captB_reg[28]  ( .D(n146), .CP(clk), .CD(n1485), .Q(captB[28]) );
  CFD2QXL \captC_reg[30]  ( .D(n116), .CP(clk), .CD(n1465), .Q(captC[30]) );
  CFD2QXL \captC_reg[28]  ( .D(n114), .CP(clk), .CD(n1466), .Q(captC[28]) );
  CFD2QXL \captA_reg[29]  ( .D(n179), .CP(clk), .CD(n1444), .Q(captA[29]) );
  CFD2QXL \captB_reg[29]  ( .D(n147), .CP(clk), .CD(n1483), .Q(captB[29]) );
  CFD2QXL \captC_reg[29]  ( .D(n115), .CP(clk), .CD(n1465), .Q(captC[29]) );
  CFD2QXL \captA_reg[27]  ( .D(n177), .CP(clk), .CD(n1445), .Q(captA[27]) );
  CFD2QXL \captB_reg[27]  ( .D(n145), .CP(clk), .CD(n1486), .Q(captB[27]) );
  CFD2QXL \captC_reg[27]  ( .D(n113), .CP(clk), .CD(n1466), .Q(captC[27]) );
  CFD2QXL \captA_reg[26]  ( .D(n176), .CP(clk), .CD(n1424), .Q(captA[26]) );
  CFD2QXL \captC_reg[26]  ( .D(n112), .CP(clk), .CD(n1467), .Q(captC[26]) );
  CFD2QXL \captB_reg[26]  ( .D(n144), .CP(clk), .CD(n1488), .Q(captB[26]) );
  CFD2QXL \captA_reg[25]  ( .D(n175), .CP(clk), .CD(n1425), .Q(captA[25]) );
  CFD2QXL \captB_reg[25]  ( .D(n143), .CP(clk), .CD(n1490), .Q(captB[25]) );
  CFD2QXL \captC_reg[25]  ( .D(n111), .CP(clk), .CD(n1467), .Q(captC[25]) );
  CFD2QXL \captA_reg[24]  ( .D(n174), .CP(clk), .CD(n1425), .Q(captA[24]) );
  CFD2QXL \captB_reg[24]  ( .D(n142), .CP(clk), .CD(n1469), .Q(captB[24]) );
  CFD2QXL \captC_reg[24]  ( .D(n110), .CP(clk), .CD(n1467), .Q(captC[24]) );
  CFD2QXL \captA_reg[23]  ( .D(n173), .CP(clk), .CD(n1426), .Q(captA[23]) );
  CFD2QXL \captB_reg[23]  ( .D(n141), .CP(clk), .CD(n1471), .Q(captB[23]) );
  CFD2QXL \captC_reg[23]  ( .D(n109), .CP(clk), .CD(n1446), .Q(captC[23]) );
  CFD2QXL \f13_reg[30]  ( .D(n1315), .CP(clk), .CD(n1480), .Q(f13[30]) );
  CFD2QXL \seen_reg[1]  ( .D(seen_d[1]), .CP(clk), .CD(n1442), .Q(stopB) );
  CFD2QXL \seen_reg[0]  ( .D(seen_d[0]), .CP(clk), .CD(n1468), .Q(stopC) );
  CFD2QXL \seen_reg[2]  ( .D(seen_d[2]), .CP(clk), .CD(n1463), .Q(stopA) );
  CFD2QXL \f34_reg[28]  ( .D(n1305), .CP(clk), .CD(n1444), .Q(f34[28]) );
  CFD2QXL \f34_reg[27]  ( .D(n1307), .CP(clk), .CD(n1445), .Q(f34[27]) );
  CFD2QXL \f34_reg[26]  ( .D(n1309), .CP(clk), .CD(n1445), .Q(f34[26]) );
  CFD2QXL \f34_reg[25]  ( .D(n1311), .CP(clk), .CD(n1424), .Q(f34[25]) );
  CFD2QXL \f34_reg[24]  ( .D(n1313), .CP(clk), .CD(n1425), .Q(f34[24]) );
  CFD2QXL \f35_reg[28]  ( .D(n1295), .CP(clk), .CD(n1484), .Q(f35[28]) );
  CFD2QXL \f35_reg[27]  ( .D(n1297), .CP(clk), .CD(n1485), .Q(f35[27]) );
  CFD2QXL \f35_reg[26]  ( .D(n1299), .CP(clk), .CD(n1487), .Q(f35[26]) );
  CFD2QXL \f35_reg[25]  ( .D(n1301), .CP(clk), .CD(n1489), .Q(f35[25]) );
  CFD2QXL \f35_reg[24]  ( .D(n1303), .CP(clk), .CD(n1468), .Q(f35[24]) );
  CFD2QXL \f44_reg[28]  ( .D(n1285), .CP(clk), .CD(n1485), .Q(f44[28]) );
  CFD2QXL \f44_reg[27]  ( .D(n1287), .CP(clk), .CD(n1486), .Q(f44[27]) );
  CFD2QXL \f44_reg[26]  ( .D(n1289), .CP(clk), .CD(n1488), .Q(f44[26]) );
  CFD2QXL \f44_reg[25]  ( .D(n1291), .CP(clk), .CD(n1489), .Q(f44[25]) );
  CFD2QXL \f44_reg[24]  ( .D(n1293), .CP(clk), .CD(n1469), .Q(f44[24]) );
  CFD2QXL \f51_reg[28]  ( .D(n1275), .CP(clk), .CD(n1484), .Q(f51[28]) );
  CFD2QXL \f51_reg[27]  ( .D(n1277), .CP(clk), .CD(n1486), .Q(f51[27]) );
  CFD2QXL \f51_reg[26]  ( .D(n1279), .CP(clk), .CD(n1487), .Q(f51[26]) );
  CFD2QXL \f51_reg[25]  ( .D(n1281), .CP(clk), .CD(n1489), .Q(f51[25]) );
  CFD2QXL \f51_reg[24]  ( .D(n1283), .CP(clk), .CD(n1468), .Q(f51[24]) );
  CFD2QXL \f62_reg[28]  ( .D(n1265), .CP(clk), .CD(n1483), .Q(f62[28]) );
  CFD2QXL \f62_reg[27]  ( .D(n1267), .CP(clk), .CD(n1485), .Q(f62[27]) );
  CFD2QXL \f62_reg[26]  ( .D(n1269), .CP(clk), .CD(n1487), .Q(f62[26]) );
  CFD2QXL \f62_reg[25]  ( .D(n1271), .CP(clk), .CD(n1488), .Q(f62[25]) );
  CFD2QXL \f62_reg[24]  ( .D(n1273), .CP(clk), .CD(n1468), .Q(f62[24]) );
  CFD2QXL \f71_reg[28]  ( .D(n1255), .CP(clk), .CD(n1484), .Q(f71[28]) );
  CFD2QXL \f71_reg[27]  ( .D(n1257), .CP(clk), .CD(n1486), .Q(f71[27]) );
  CFD2QXL \f71_reg[26]  ( .D(n1259), .CP(clk), .CD(n1487), .Q(f71[26]) );
  CFD2QXL \f34_reg[9]  ( .D(n1261), .CP(clk), .CD(n1457), .Q(f34[9]) );
  CFD2QXL \f34_reg[11]  ( .D(n1263), .CP(clk), .CD(n1434), .Q(f34[11]) );
  CFD2QXL \f34_reg[0]  ( .D(n1245), .CP(clk), .CD(n1463), .Q(f34[0]) );
  CFD2QXL \f35_reg[0]  ( .D(n1247), .CP(clk), .CD(n1441), .Q(f35[0]) );
  CFD2QXL \f44_reg[0]  ( .D(n1249), .CP(clk), .CD(n1441), .Q(f44[0]) );
  CFD2QXL \f51_reg[0]  ( .D(n1251), .CP(clk), .CD(n1441), .Q(f51[0]) );
  CFD2QXL \f62_reg[0]  ( .D(n1253), .CP(clk), .CD(n1440), .Q(f62[0]) );
  CFD2QXL \f34_reg[3]  ( .D(n1235), .CP(clk), .CD(n1461), .Q(f34[3]) );
  CFD2QXL \f35_reg[11]  ( .D(n1237), .CP(clk), .CD(n1490), .Q(f35[11]) );
  CFD2QXL \f44_reg[11]  ( .D(n1239), .CP(clk), .CD(n1491), .Q(f44[11]) );
  CFD2QXL \f51_reg[11]  ( .D(n1241), .CP(clk), .CD(n1490), .Q(f51[11]) );
  CFD2QXL \f62_reg[11]  ( .D(n1243), .CP(clk), .CD(n1510), .Q(f62[11]) );
  CFD2QXL \f35_reg[9]  ( .D(n1225), .CP(clk), .CD(n1493), .Q(f35[9]) );
  CFD2QXL \f44_reg[9]  ( .D(n1227), .CP(clk), .CD(n1494), .Q(f44[9]) );
  CFD2QXL \f51_reg[9]  ( .D(n1229), .CP(clk), .CD(n1493), .Q(f51[9]) );
  CFD2QXL \f62_reg[9]  ( .D(n1231), .CP(clk), .CD(n1493), .Q(f62[9]) );
  CFD2QXL \f35_reg[3]  ( .D(n1233), .CP(clk), .CD(n1436), .Q(f35[3]) );
  CFD2QXL \f44_reg[3]  ( .D(n1215), .CP(clk), .CD(n1437), .Q(f44[3]) );
  CFD2QXL \f51_reg[3]  ( .D(n1217), .CP(clk), .CD(n1436), .Q(f51[3]) );
  CFD2QXL \f62_reg[3]  ( .D(n1219), .CP(clk), .CD(n1436), .Q(f62[3]) );
  CFD2QXL \f34_reg[1]  ( .D(n1221), .CP(clk), .CD(n1462), .Q(f34[1]) );
  CFD2QXL \f71_reg[3]  ( .D(n1223), .CP(clk), .CD(n1436), .Q(f71[3]) );
  CFD2QXL \f71_reg[1]  ( .D(n1205), .CP(clk), .CD(n1439), .Q(f71[1]) );
  CFD2QXL \f34_reg[23]  ( .D(n1207), .CP(clk), .CD(n1426), .Q(f34[23]) );
  CFD2QXL \f34_reg[21]  ( .D(n1209), .CP(clk), .CD(n1427), .Q(f34[21]) );
  CFD2QXL \f34_reg[19]  ( .D(n1211), .CP(clk), .CD(n1428), .Q(f34[19]) );
  CFD2QXL \f34_reg[17]  ( .D(n1213), .CP(clk), .CD(n1430), .Q(f34[17]) );
  CFD2QXL \f34_reg[16]  ( .D(n1195), .CP(clk), .CD(n1430), .Q(f34[16]) );
  CFD2QXL \f34_reg[15]  ( .D(n1197), .CP(clk), .CD(n1431), .Q(f34[15]) );
  CFD2QXL \f34_reg[14]  ( .D(n1199), .CP(clk), .CD(n1432), .Q(f34[14]) );
  CFD2QXL \f34_reg[13]  ( .D(n1201), .CP(clk), .CD(n1432), .Q(f34[13]) );
  CFD2QXL \f34_reg[12]  ( .D(n1203), .CP(clk), .CD(n1433), .Q(f34[12]) );
  CFD2QXL \f34_reg[8]  ( .D(n1185), .CP(clk), .CD(n1458), .Q(f34[8]) );
  CFD2QXL \f34_reg[7]  ( .D(n1187), .CP(clk), .CD(n1458), .Q(f34[7]) );
  CFD2QXL \f34_reg[5]  ( .D(n1189), .CP(clk), .CD(n1459), .Q(f34[5]) );
  CFD2QXL \f34_reg[4]  ( .D(n1191), .CP(clk), .CD(n1460), .Q(f34[4]) );
  CFD2QXL \f35_reg[23]  ( .D(n1193), .CP(clk), .CD(n1470), .Q(f35[23]) );
  CFD2QXL \f35_reg[21]  ( .D(n1175), .CP(clk), .CD(n1473), .Q(f35[21]) );
  CFD2QXL \f35_reg[19]  ( .D(n1177), .CP(clk), .CD(n1476), .Q(f35[19]) );
  CFD2QXL \f35_reg[17]  ( .D(n1179), .CP(clk), .CD(n1501), .Q(f35[17]) );
  CFD2QXL \f35_reg[16]  ( .D(n1181), .CP(clk), .CD(n1503), .Q(f35[16]) );
  CFD2QXL \f35_reg[8]  ( .D(n1183), .CP(clk), .CD(n1495), .Q(f35[8]) );
  CFD2QXL \f35_reg[5]  ( .D(n1165), .CP(clk), .CD(n1499), .Q(f35[5]) );
  CFD2QXL \f35_reg[4]  ( .D(n1167), .CP(clk), .CD(n1440), .Q(f35[4]) );
  CFD2QXL \f44_reg[23]  ( .D(n1169), .CP(clk), .CD(n1470), .Q(f44[23]) );
  CFD2QXL \f44_reg[21]  ( .D(n1171), .CP(clk), .CD(n1474), .Q(f44[21]) );
  CFD2QXL \f44_reg[19]  ( .D(n1173), .CP(clk), .CD(n1477), .Q(f44[19]) );
  CFD2QXL \f44_reg[17]  ( .D(n1155), .CP(clk), .CD(n1502), .Q(f44[17]) );
  CFD2QXL \f44_reg[16]  ( .D(n1157), .CP(clk), .CD(n1503), .Q(f44[16]) );
  CFD2QXL \f44_reg[8]  ( .D(n1159), .CP(clk), .CD(n1495), .Q(f44[8]) );
  CFD2QXL \f44_reg[5]  ( .D(n1161), .CP(clk), .CD(n1500), .Q(f44[5]) );
  CFD2QXL \f44_reg[4]  ( .D(n1163), .CP(clk), .CD(n1435), .Q(f44[4]) );
  CFD2QXL \f51_reg[23]  ( .D(n1145), .CP(clk), .CD(n1470), .Q(f51[23]) );
  CFD2QXL \f51_reg[21]  ( .D(n1147), .CP(clk), .CD(n1473), .Q(f51[21]) );
  CFD2QXL \f51_reg[19]  ( .D(n1149), .CP(clk), .CD(n1476), .Q(f51[19]) );
  CFD2QXL \f51_reg[17]  ( .D(n1151), .CP(clk), .CD(n1502), .Q(f51[17]) );
  CFD2QXL \f51_reg[16]  ( .D(n1153), .CP(clk), .CD(n1503), .Q(f51[16]) );
  CFD2QXL \f51_reg[8]  ( .D(n1135), .CP(clk), .CD(n1495), .Q(f51[8]) );
  CFD2QXL \f51_reg[5]  ( .D(n1137), .CP(clk), .CD(n1500), .Q(f51[5]) );
  CFD2QXL \f51_reg[4]  ( .D(n1139), .CP(clk), .CD(n1435), .Q(f51[4]) );
  CFD2QXL \f62_reg[23]  ( .D(n1141), .CP(clk), .CD(n1469), .Q(f62[23]) );
  CFD2QXL \f62_reg[21]  ( .D(n1143), .CP(clk), .CD(n1472), .Q(f62[21]) );
  CFD2QXL \f62_reg[19]  ( .D(n1125), .CP(clk), .CD(n1476), .Q(f62[19]) );
  CFD2QXL \f62_reg[17]  ( .D(n1127), .CP(clk), .CD(n1501), .Q(f62[17]) );
  CFD2QXL \f62_reg[16]  ( .D(n1129), .CP(clk), .CD(n1502), .Q(f62[16]) );
  CFD2QXL \f62_reg[8]  ( .D(n1131), .CP(clk), .CD(n1494), .Q(f62[8]) );
  CFD2QXL \f62_reg[5]  ( .D(n1133), .CP(clk), .CD(n1499), .Q(f62[5]) );
  CFD2QXL \f62_reg[4]  ( .D(n1115), .CP(clk), .CD(n1501), .Q(f62[4]) );
  CFD2QXL \f71_reg[25]  ( .D(n1117), .CP(clk), .CD(n1489), .Q(f71[25]) );
  CFD2QXL \f71_reg[24]  ( .D(n1119), .CP(clk), .CD(n1468), .Q(f71[24]) );
  CFD2QXL \f71_reg[23]  ( .D(n1121), .CP(clk), .CD(n1470), .Q(f71[23]) );
  CFD2QXL \f71_reg[21]  ( .D(n1123), .CP(clk), .CD(n1473), .Q(f71[21]) );
  CFD2QXL \f71_reg[20]  ( .D(n1105), .CP(clk), .CD(n1475), .Q(f71[20]) );
  CFD2QXL \f71_reg[19]  ( .D(n1107), .CP(clk), .CD(n1476), .Q(f71[19]) );
  CFD2QXL \f71_reg[17]  ( .D(n1109), .CP(clk), .CD(n1501), .Q(f71[17]) );
  CFD2QXL \f71_reg[16]  ( .D(n1111), .CP(clk), .CD(n1503), .Q(f71[16]) );
  CFD2QXL \f71_reg[15]  ( .D(n1113), .CP(clk), .CD(n1504), .Q(f71[15]) );
  CFD2QXL \f71_reg[14]  ( .D(n1095), .CP(clk), .CD(n1506), .Q(f71[14]) );
  CFD2QXL \f71_reg[13]  ( .D(n1097), .CP(clk), .CD(n1508), .Q(f71[13]) );
  CFD2QXL \f71_reg[12]  ( .D(n1099), .CP(clk), .CD(n1510), .Q(f71[12]) );
  CFD2QXL \f71_reg[11]  ( .D(n1101), .CP(clk), .CD(n1490), .Q(f71[11]) );
  CFD2QXL \f71_reg[10]  ( .D(n1103), .CP(clk), .CD(n1492), .Q(f71[10]) );
  CFD2QXL \f71_reg[9]  ( .D(n1085), .CP(clk), .CD(n1493), .Q(f71[9]) );
  CFD2QXL \f71_reg[8]  ( .D(n1087), .CP(clk), .CD(n1495), .Q(f71[8]) );
  CFD2QXL \f71_reg[7]  ( .D(n1089), .CP(clk), .CD(n1496), .Q(f71[7]) );
  CFD2QXL \f71_reg[4]  ( .D(n1091), .CP(clk), .CD(n1435), .Q(f71[4]) );
  CFD2QXL \f71_reg[0]  ( .D(n1093), .CP(clk), .CD(n1441), .Q(f71[0]) );
  CFD2QXL \f35_reg[10]  ( .D(n1075), .CP(clk), .CD(n1491), .Q(f35[10]) );
  CFD2QXL \f44_reg[10]  ( .D(n1077), .CP(clk), .CD(n1492), .Q(f44[10]) );
  CFD2QXL \f51_reg[10]  ( .D(n1079), .CP(clk), .CD(n1492), .Q(f51[10]) );
  CFD2QXL \f62_reg[10]  ( .D(n1081), .CP(clk), .CD(n1491), .Q(f62[10]) );
  CFD2QXL \f35_reg[15]  ( .D(n1083), .CP(clk), .CD(n1504), .Q(f35[15]) );
  CFD2QXL \f44_reg[15]  ( .D(n1065), .CP(clk), .CD(n1505), .Q(f44[15]) );
  CFD2QXL \f51_reg[15]  ( .D(n1067), .CP(clk), .CD(n1504), .Q(f51[15]) );
  CFD2QXL \f62_reg[15]  ( .D(n1069), .CP(clk), .CD(n1504), .Q(f62[15]) );
  CFD2QXL \f35_reg[13]  ( .D(n1071), .CP(clk), .CD(n1507), .Q(f35[13]) );
  CFD2QXL \f44_reg[13]  ( .D(n1073), .CP(clk), .CD(n1509), .Q(f44[13]) );
  CFD2QXL \f51_reg[13]  ( .D(n1055), .CP(clk), .CD(n1508), .Q(f51[13]) );
  CFD2QXL \f62_reg[13]  ( .D(n1057), .CP(clk), .CD(n1507), .Q(f62[13]) );
  CFD2QXL \f35_reg[7]  ( .D(n1059), .CP(clk), .CD(n1496), .Q(f35[7]) );
  CFD2QXL \f44_reg[7]  ( .D(n1061), .CP(clk), .CD(n1497), .Q(f44[7]) );
  CFD2QXL \f51_reg[7]  ( .D(n1063), .CP(clk), .CD(n1496), .Q(f51[7]) );
  CFD2QXL \f62_reg[7]  ( .D(n1045), .CP(clk), .CD(n1496), .Q(f62[7]) );
  CFD2QXL \f35_reg[14]  ( .D(n1047), .CP(clk), .CD(n1506), .Q(f35[14]) );
  CFD2QXL \f44_reg[14]  ( .D(n1049), .CP(clk), .CD(n1507), .Q(f44[14]) );
  CFD2QXL \f51_reg[14]  ( .D(n1051), .CP(clk), .CD(n1506), .Q(f51[14]) );
  CFD2QXL \f62_reg[14]  ( .D(n1053), .CP(clk), .CD(n1505), .Q(f62[14]) );
  CFD2QXL \f35_reg[12]  ( .D(n1035), .CP(clk), .CD(n1510), .Q(f35[12]) );
  CFD2QXL \f44_reg[12]  ( .D(n1037), .CP(clk), .CD(n1510), .Q(f44[12]) );
  CFD2QXL \f51_reg[12]  ( .D(n1039), .CP(clk), .CD(n1510), .Q(f51[12]) );
  CFD2QXL \f62_reg[12]  ( .D(n1041), .CP(clk), .CD(n1508), .Q(f62[12]) );
  CFD2QXL \f34_reg[10]  ( .D(n1043), .CP(clk), .CD(n1434), .Q(f34[10]) );
  CFD2QXL \f35_reg[1]  ( .D(n1025), .CP(clk), .CD(n1439), .Q(f35[1]) );
  CFD2QXL \f51_reg[1]  ( .D(n1027), .CP(clk), .CD(n1439), .Q(f51[1]) );
  CFD2QXL \f62_reg[1]  ( .D(n1029), .CP(clk), .CD(n1439), .Q(f62[1]) );
  CFD2QXL \f34_reg[22]  ( .D(n1031), .CP(clk), .CD(n1426), .Q(f34[22]) );
  CFD2QXL \f34_reg[20]  ( .D(n1033), .CP(clk), .CD(n1428), .Q(f34[20]) );
  CFD2QXL \f34_reg[18]  ( .D(n1015), .CP(clk), .CD(n1429), .Q(f34[18]) );
  CFD2QXL \f34_reg[6]  ( .D(n1017), .CP(clk), .CD(n1459), .Q(f34[6]) );
  CFD2QXL \f34_reg[2]  ( .D(n1019), .CP(clk), .CD(n1461), .Q(f34[2]) );
  CFD2QXL \f35_reg[22]  ( .D(n1021), .CP(clk), .CD(n1471), .Q(f35[22]) );
  CFD2QXL \f35_reg[20]  ( .D(n1023), .CP(clk), .CD(n1474), .Q(f35[20]) );
  CFD2QXL \f35_reg[18]  ( .D(n1005), .CP(clk), .CD(n1478), .Q(f35[18]) );
  CFD2QXL \f35_reg[6]  ( .D(n1007), .CP(clk), .CD(n1498), .Q(f35[6]) );
  CFD2QXL \f35_reg[2]  ( .D(n1009), .CP(clk), .CD(n1438), .Q(f35[2]) );
  CFD2QXL \f44_reg[22]  ( .D(n1011), .CP(clk), .CD(n1472), .Q(f44[22]) );
  CFD2QXL \f44_reg[20]  ( .D(n1013), .CP(clk), .CD(n1475), .Q(f44[20]) );
  CFD2QXL \f44_reg[18]  ( .D(n995), .CP(clk), .CD(n1478), .Q(f44[18]) );
  CFD2QXL \f44_reg[6]  ( .D(n997), .CP(clk), .CD(n1498), .Q(f44[6]) );
  CFD2QXL \f44_reg[2]  ( .D(n999), .CP(clk), .CD(n1438), .Q(f44[2]) );
  CFD2QXL \f51_reg[22]  ( .D(n1001), .CP(clk), .CD(n1472), .Q(f51[22]) );
  CFD2QXL \f51_reg[20]  ( .D(n1003), .CP(clk), .CD(n1475), .Q(f51[20]) );
  CFD2QXL \f51_reg[18]  ( .D(n985), .CP(clk), .CD(n1478), .Q(f51[18]) );
  CFD2QXL \f51_reg[6]  ( .D(n987), .CP(clk), .CD(n1498), .Q(f51[6]) );
  CFD2QXL \f51_reg[2]  ( .D(n989), .CP(clk), .CD(n1438), .Q(f51[2]) );
  CFD2QXL \f62_reg[22]  ( .D(n991), .CP(clk), .CD(n1471), .Q(f62[22]) );
  CFD2QXL \f62_reg[20]  ( .D(n993), .CP(clk), .CD(n1474), .Q(f62[20]) );
  CFD2QXL \f62_reg[18]  ( .D(n975), .CP(clk), .CD(n1477), .Q(f62[18]) );
  CFD2QXL \f62_reg[6]  ( .D(n977), .CP(clk), .CD(n1497), .Q(f62[6]) );
  CFD2QXL \f62_reg[2]  ( .D(n979), .CP(clk), .CD(n1437), .Q(f62[2]) );
  CFD2QXL \f71_reg[22]  ( .D(n981), .CP(clk), .CD(n1471), .Q(f71[22]) );
  CFD2QXL \f71_reg[18]  ( .D(n983), .CP(clk), .CD(n1478), .Q(f71[18]) );
  CFD2QXL \f71_reg[6]  ( .D(n964), .CP(clk), .CD(n1498), .Q(f71[6]) );
  CFD2QXL \f71_reg[5]  ( .D(n966), .CP(clk), .CD(n1500), .Q(f71[5]) );
  CFD2QXL \f71_reg[2]  ( .D(n968), .CP(clk), .CD(n1438), .Q(f71[2]) );
  CFD2QXL \f13_reg[14]  ( .D(n970), .CP(clk), .CD(n1506), .Q(f13[14]) );
  CFD2QXL \f13_reg[13]  ( .D(n972), .CP(clk), .CD(n1508), .Q(f13[13]) );
  CFD2QXL \f13_reg[10]  ( .D(n957), .CP(clk), .CD(n1491), .Q(f13[10]) );
  CFD2QXL \f13_reg[5]  ( .D(n959), .CP(clk), .CD(n1499), .Q(f13[5]) );
  CFD2QXL \f13_reg[4]  ( .D(n962), .CP(clk), .CD(n1446), .Q(f13[4]) );
  CFD2QXL \f13_reg[2]  ( .D(n955), .CP(clk), .CD(n1438), .Q(f13[2]) );
  CFD2QXL \f14_reg[27]  ( .D(w2[27]), .CP(clk), .CD(n1488), .Q(f14[27]) );
  CFD2QXL \f36_reg[15]  ( .D(n951), .CP(clk), .CD(n1431), .Q(f36[15]) );
  CFD2QXL \f36_reg[14]  ( .D(n953), .CP(clk), .CD(n1431), .Q(f36[14]) );
  CFD2QXL \f36_reg[10]  ( .D(n943), .CP(clk), .CD(n1434), .Q(f36[10]) );
  CFD2QXL \f36_reg[11]  ( .D(n945), .CP(clk), .CD(n1433), .Q(f36[11]) );
  CFD2QXL \f36_reg[6]  ( .D(n941), .CP(clk), .CD(n1459), .Q(f36[6]) );
  CFD2QXL \f32_reg[28]  ( .D(w8[28]), .CP(clk), .CD(n1484), .Q(f32[28]) );
  CFD2QXL \f32_reg[27]  ( .D(w8[27]), .CP(clk), .CD(n1485), .Q(f32[27]) );
  CFD2QXL \f32_reg[26]  ( .D(w8[26]), .CP(clk), .CD(n1487), .Q(f32[26]) );
  CFD2QXL \f32_reg[25]  ( .D(w8[25]), .CP(clk), .CD(n1489), .Q(f32[25]) );
  CFD2QXL \f32_reg[24]  ( .D(w8[24]), .CP(clk), .CD(n1468), .Q(f32[24]) );
  CFD2QXL \f46_reg[28]  ( .D(n939), .CP(clk), .CD(n1466), .Q(f46[28]) );
  CFD2QXL \f46_reg[27]  ( .D(n931), .CP(clk), .CD(n1466), .Q(f46[27]) );
  CFD2QXL \f46_reg[26]  ( .D(n933), .CP(clk), .CD(n1467), .Q(f46[26]) );
  CFD2QXL \f46_reg[25]  ( .D(n935), .CP(clk), .CD(n1467), .Q(f46[25]) );
  CFD2QXL \f46_reg[24]  ( .D(n937), .CP(clk), .CD(n1446), .Q(f46[24]) );
  CFD2QXL \f53_reg[28]  ( .D(w11[28]), .CP(clk), .CD(n1444), .Q(f53[28]) );
  CFD2QXL \f53_reg[27]  ( .D(w11[27]), .CP(clk), .CD(n1444), .Q(f53[27]) );
  CFD2QXL \f53_reg[26]  ( .D(w11[26]), .CP(clk), .CD(n1445), .Q(f53[26]) );
  CFD2QXL \f53_reg[25]  ( .D(w11[25]), .CP(clk), .CD(n1424), .Q(f53[25]) );
  CFD2QXL \f53_reg[24]  ( .D(w11[24]), .CP(clk), .CD(n1425), .Q(f53[24]) );
  CFD2QXL \f63_reg[28]  ( .D(n929), .CP(clk), .CD(n1484), .Q(f63[28]) );
  CFD2QXL \f63_reg[27]  ( .D(n921), .CP(clk), .CD(n1486), .Q(f63[27]) );
  CFD2QXL \f63_reg[26]  ( .D(n923), .CP(clk), .CD(n1488), .Q(f63[26]) );
  CFD2QXL \f63_reg[25]  ( .D(n925), .CP(clk), .CD(n1489), .Q(f63[25]) );
  CFD2QXL \f63_reg[24]  ( .D(n927), .CP(clk), .CD(n1469), .Q(f63[24]) );
  CFD2QXL \f72_reg[28]  ( .D(s72[28]), .CP(clk), .CD(n1483), .Q(f72[28]) );
  CFD2QXL \f72_reg[27]  ( .D(s72[27]), .CP(clk), .CD(n1485), .Q(f72[27]) );
  CFD2QXL \f72_reg[26]  ( .D(s72[26]), .CP(clk), .CD(n1487), .Q(f72[26]) );
  CFD2QXL \f32_reg[1]  ( .D(w8[1]), .CP(clk), .CD(n1439), .Q(f32[1]) );
  CFD2QXL \f53_reg[1]  ( .D(w11[1]), .CP(clk), .CD(n1462), .Q(f53[1]) );
  CFD2QXL \f63_reg[1]  ( .D(n919), .CP(clk), .CD(n1440), .Q(f63[1]) );
  CFD2QXL \f32_reg[7]  ( .D(w8[7]), .CP(clk), .CD(n1496), .Q(f32[7]) );
  CFD2QXL \f46_reg[7]  ( .D(n915), .CP(clk), .CD(n1453), .Q(f46[7]) );
  CFD2QXL \f53_reg[7]  ( .D(w11[7]), .CP(clk), .CD(n1458), .Q(f53[7]) );
  CFD2QXL \f63_reg[7]  ( .D(n917), .CP(clk), .CD(n1497), .Q(f63[7]) );
  CFD2QXL \f32_reg[13]  ( .D(w8[13]), .CP(clk), .CD(n1507), .Q(f32[13]) );
  CFD2QXL \f46_reg[13]  ( .D(n909), .CP(clk), .CD(n1451), .Q(f46[13]) );
  CFD2QXL \f53_reg[13]  ( .D(w11[13]), .CP(clk), .CD(n1432), .Q(f53[13]) );
  CFD2QXL \f63_reg[13]  ( .D(n911), .CP(clk), .CD(n1508), .Q(f63[13]) );
  CFD2QXL \f32_reg[15]  ( .D(w8[15]), .CP(clk), .CD(n1504), .Q(f32[15]) );
  CFD2QXL \f46_reg[15]  ( .D(n913), .CP(clk), .CD(n1450), .Q(f46[15]) );
  CFD2QXL \f53_reg[15]  ( .D(w11[15]), .CP(clk), .CD(n1431), .Q(f53[15]) );
  CFD2QXL \f63_reg[15]  ( .D(n905), .CP(clk), .CD(n1505), .Q(f63[15]) );
  CFD2QXL \f32_reg[0]  ( .D(w8[0]), .CP(clk), .CD(n1441), .Q(f32[0]) );
  CFD2QXL \f46_reg[0]  ( .D(n907), .CP(clk), .CD(n1456), .Q(f46[0]) );
  CFD2QXL \f53_reg[0]  ( .D(w11[0]), .CP(clk), .CD(n1463), .Q(f53[0]) );
  CFD2QXL \f63_reg[0]  ( .D(n899), .CP(clk), .CD(n1441), .Q(f63[0]) );
  CFD2QXL \f32_reg[3]  ( .D(w8[3]), .CP(clk), .CD(n1436), .Q(f32[3]) );
  CFD2QXL \f46_reg[3]  ( .D(n901), .CP(clk), .CD(n1455), .Q(f46[3]) );
  CFD2QXL \f53_reg[3]  ( .D(w11[3]), .CP(clk), .CD(n1460), .Q(f53[3]) );
  CFD2QXL \f63_reg[3]  ( .D(n903), .CP(clk), .CD(n1437), .Q(f63[3]) );
  CFD2QXL \f32_reg[11]  ( .D(w8[11]), .CP(clk), .CD(n1495), .Q(f32[11]) );
  CFD2QXL \f46_reg[11]  ( .D(n895), .CP(clk), .CD(n1452), .Q(f46[11]) );
  CFD2QXL \f53_reg[11]  ( .D(w11[11]), .CP(clk), .CD(n1433), .Q(f53[11]) );
  CFD2QXL \f63_reg[11]  ( .D(n897), .CP(clk), .CD(n1490), .Q(f63[11]) );
  CFD2QXL \f72_reg[3]  ( .D(s72[3]), .CP(clk), .CD(n1436), .Q(f72[3]) );
  CFD2QXL \f72_reg[1]  ( .D(s72[1]), .CP(clk), .CD(n1439), .Q(f72[1]) );
  CFD2QXL \f32_reg[23]  ( .D(w8[23]), .CP(clk), .CD(n1470), .Q(f32[23]) );
  CFD2QXL \f32_reg[21]  ( .D(w8[21]), .CP(clk), .CD(n1473), .Q(f32[21]) );
  CFD2QXL \f32_reg[19]  ( .D(w8[19]), .CP(clk), .CD(n1476), .Q(f32[19]) );
  CFD2QXL \f32_reg[17]  ( .D(w8[17]), .CP(clk), .CD(n1501), .Q(f32[17]) );
  CFD2QXL \f32_reg[16]  ( .D(w8[16]), .CP(clk), .CD(n1503), .Q(f32[16]) );
  CFD2QXL \f32_reg[8]  ( .D(w8[8]), .CP(clk), .CD(n1494), .Q(f32[8]) );
  CFD2QXL \f32_reg[5]  ( .D(w8[5]), .CP(clk), .CD(n1499), .Q(f32[5]) );
  CFD2QXL \f32_reg[4]  ( .D(w8[4]), .CP(clk), .CD(n1501), .Q(f32[4]) );
  CFD2QXL \f46_reg[23]  ( .D(n893), .CP(clk), .CD(n1446), .Q(f46[23]) );
  CFD2QXL \f46_reg[21]  ( .D(n883), .CP(clk), .CD(n1447), .Q(f46[21]) );
  CFD2QXL \f46_reg[19]  ( .D(n885), .CP(clk), .CD(n1448), .Q(f46[19]) );
  CFD2QXL \f46_reg[17]  ( .D(n887), .CP(clk), .CD(n1449), .Q(f46[17]) );
  CFD2QXL \f46_reg[16]  ( .D(n889), .CP(clk), .CD(n1449), .Q(f46[16]) );
  CFD2QXL \f46_reg[8]  ( .D(n891), .CP(clk), .CD(n1453), .Q(f46[8]) );
  CFD2QXL \f46_reg[5]  ( .D(n879), .CP(clk), .CD(n1454), .Q(f46[5]) );
  CFD2QXL \f46_reg[4]  ( .D(n881), .CP(clk), .CD(n1455), .Q(f46[4]) );
  CFD2QXL \f53_reg[23]  ( .D(w11[23]), .CP(clk), .CD(n1426), .Q(f53[23]) );
  CFD2QXL \f53_reg[21]  ( .D(w11[21]), .CP(clk), .CD(n1427), .Q(f53[21]) );
  CFD2QXL \f53_reg[19]  ( .D(w11[19]), .CP(clk), .CD(n1428), .Q(f53[19]) );
  CFD2QXL \f53_reg[17]  ( .D(w11[17]), .CP(clk), .CD(n1429), .Q(f53[17]) );
  CFD2QXL \f53_reg[16]  ( .D(w11[16]), .CP(clk), .CD(n1430), .Q(f53[16]) );
  CFD2QXL \f53_reg[8]  ( .D(w11[8]), .CP(clk), .CD(n1457), .Q(f53[8]) );
  CFD2QXL \f53_reg[5]  ( .D(w11[5]), .CP(clk), .CD(n1459), .Q(f53[5]) );
  CFD2QXL \f53_reg[4]  ( .D(w11[4]), .CP(clk), .CD(n1460), .Q(f53[4]) );
  CFD2QXL \f63_reg[23]  ( .D(n869), .CP(clk), .CD(n1470), .Q(f63[23]) );
  CFD2QXL \f63_reg[21]  ( .D(n871), .CP(clk), .CD(n1473), .Q(f63[21]) );
  CFD2QXL \f63_reg[19]  ( .D(n873), .CP(clk), .CD(n1477), .Q(f63[19]) );
  CFD2QXL \f63_reg[17]  ( .D(n875), .CP(clk), .CD(n1502), .Q(f63[17]) );
  CFD2QXL \f63_reg[16]  ( .D(n877), .CP(clk), .CD(n1503), .Q(f63[16]) );
  CFD2QXL \f63_reg[8]  ( .D(n863), .CP(clk), .CD(n1495), .Q(f63[8]) );
  CFD2QXL \f63_reg[5]  ( .D(n865), .CP(clk), .CD(n1500), .Q(f63[5]) );
  CFD2QXL \f63_reg[4]  ( .D(n867), .CP(clk), .CD(n1435), .Q(f63[4]) );
  CFD2QXL \f72_reg[25]  ( .D(s72[25]), .CP(clk), .CD(n1488), .Q(f72[25]) );
  CFD2QXL \f72_reg[24]  ( .D(s72[24]), .CP(clk), .CD(n1468), .Q(f72[24]) );
  CFD2QXL \f72_reg[23]  ( .D(s72[23]), .CP(clk), .CD(n1469), .Q(f72[23]) );
  CFD2QXL \f72_reg[21]  ( .D(s72[21]), .CP(clk), .CD(n1472), .Q(f72[21]) );
  CFD2QXL \f72_reg[20]  ( .D(s72[20]), .CP(clk), .CD(n1474), .Q(f72[20]) );
  CFD2QXL \f72_reg[19]  ( .D(s72[19]), .CP(clk), .CD(n1476), .Q(f72[19]) );
  CFD2QXL \f72_reg[17]  ( .D(s72[17]), .CP(clk), .CD(n1506), .Q(f72[17]) );
  CFD2QXL \f72_reg[16]  ( .D(s72[16]), .CP(clk), .CD(n1502), .Q(f72[16]) );
  CFD2QXL \f72_reg[15]  ( .D(s72[15]), .CP(clk), .CD(n1504), .Q(f72[15]) );
  CFD2QXL \f72_reg[14]  ( .D(s72[14]), .CP(clk), .CD(n1505), .Q(f72[14]) );
  CFD2QXL \f72_reg[13]  ( .D(s72[13]), .CP(clk), .CD(n1507), .Q(f72[13]) );
  CFD2QXL \f72_reg[12]  ( .D(s72[12]), .CP(clk), .CD(n1509), .Q(f72[12]) );
  CFD2QXL \f72_reg[11]  ( .D(s72[11]), .CP(clk), .CD(n1510), .Q(f72[11]) );
  CFD2QXL \f72_reg[10]  ( .D(s72[10]), .CP(clk), .CD(n1491), .Q(f72[10]) );
  CFD2QXL \f72_reg[9]  ( .D(s72[9]), .CP(clk), .CD(n1493), .Q(f72[9]) );
  CFD2QXL \f72_reg[8]  ( .D(s72[8]), .CP(clk), .CD(n1494), .Q(f72[8]) );
  CFD2QXL \f72_reg[7]  ( .D(s72[7]), .CP(clk), .CD(n1496), .Q(f72[7]) );
  CFD2QXL \f72_reg[4]  ( .D(s72[4]), .CP(clk), .CD(n1501), .Q(f72[4]) );
  CFD2QXL \f72_reg[0]  ( .D(s72[0]), .CP(clk), .CD(n1440), .Q(f72[0]) );
  CFD2QXL \f32_reg[10]  ( .D(w8[10]), .CP(clk), .CD(n1491), .Q(f32[10]) );
  CFD2QXL \f46_reg[10]  ( .D(n861), .CP(clk), .CD(n1452), .Q(f46[10]) );
  CFD2QXL \f53_reg[10]  ( .D(w11[10]), .CP(clk), .CD(n1434), .Q(f53[10]) );
  CFD2QXL \f63_reg[10]  ( .D(n855), .CP(clk), .CD(n1492), .Q(f63[10]) );
  CFD2QXL \f32_reg[14]  ( .D(w8[14]), .CP(clk), .CD(n1506), .Q(f32[14]) );
  CFD2QXL \f46_reg[14]  ( .D(n857), .CP(clk), .CD(n1450), .Q(f46[14]) );
  CFD2QXL \f53_reg[14]  ( .D(w11[14]), .CP(clk), .CD(n1431), .Q(f53[14]) );
  CFD2QXL \f63_reg[14]  ( .D(n859), .CP(clk), .CD(n1506), .Q(f63[14]) );
  CFD2QXL \f32_reg[12]  ( .D(w8[12]), .CP(clk), .CD(n1509), .Q(f32[12]) );
  CFD2QXL \f46_reg[12]  ( .D(n851), .CP(clk), .CD(n1451), .Q(f46[12]) );
  CFD2QXL \f53_reg[12]  ( .D(w11[12]), .CP(clk), .CD(n1433), .Q(f53[12]) );
  CFD2QXL \f63_reg[12]  ( .D(n853), .CP(clk), .CD(n1509), .Q(f63[12]) );
  CFD2QXL \f32_reg[22]  ( .D(w8[22]), .CP(clk), .CD(n1471), .Q(f32[22]) );
  CFD2QXL \f32_reg[20]  ( .D(w8[20]), .CP(clk), .CD(n1474), .Q(f32[20]) );
  CFD2QXL \f32_reg[18]  ( .D(w8[18]), .CP(clk), .CD(n1477), .Q(f32[18]) );
  CFD2QXL \f32_reg[6]  ( .D(w8[6]), .CP(clk), .CD(n1498), .Q(f32[6]) );
  CFD2QXL \f32_reg[2]  ( .D(w8[2]), .CP(clk), .CD(n1437), .Q(f32[2]) );
  CFD2QXL \f46_reg[22]  ( .D(n849), .CP(clk), .CD(n1447), .Q(f46[22]) );
  CFD2QXL \f46_reg[20]  ( .D(n841), .CP(clk), .CD(n1447), .Q(f46[20]) );
  CFD2QXL \f46_reg[18]  ( .D(n843), .CP(clk), .CD(n1448), .Q(f46[18]) );
  CFD2QXL \f46_reg[6]  ( .D(n845), .CP(clk), .CD(n1454), .Q(f46[6]) );
  CFD2QXL \f46_reg[2]  ( .D(n847), .CP(clk), .CD(n1456), .Q(f46[2]) );
  CFD2QXL \f53_reg[22]  ( .D(w11[22]), .CP(clk), .CD(n1426), .Q(f53[22]) );
  CFD2QXL \f53_reg[20]  ( .D(w11[20]), .CP(clk), .CD(n1427), .Q(f53[20]) );
  CFD2QXL \f53_reg[18]  ( .D(w11[18]), .CP(clk), .CD(n1429), .Q(f53[18]) );
  CFD2QXL \f53_reg[6]  ( .D(w11[6]), .CP(clk), .CD(n1459), .Q(f53[6]) );
  CFD2QXL \f53_reg[2]  ( .D(w11[2]), .CP(clk), .CD(n1461), .Q(f53[2]) );
  CFD2QXL \f63_reg[22]  ( .D(n839), .CP(clk), .CD(n1472), .Q(f63[22]) );
  CFD2QXL \f63_reg[20]  ( .D(n831), .CP(clk), .CD(n1475), .Q(f63[20]) );
  CFD2QXL \f63_reg[18]  ( .D(n833), .CP(clk), .CD(n1478), .Q(f63[18]) );
  CFD2QXL \f63_reg[6]  ( .D(n835), .CP(clk), .CD(n1498), .Q(f63[6]) );
  CFD2QXL \f63_reg[2]  ( .D(n837), .CP(clk), .CD(n1438), .Q(f63[2]) );
  CFD2QXL \f72_reg[22]  ( .D(s72[22]), .CP(clk), .CD(n1471), .Q(f72[22]) );
  CFD2QXL \f72_reg[18]  ( .D(s72[18]), .CP(clk), .CD(n1477), .Q(f72[18]) );
  CFD2QXL \f72_reg[6]  ( .D(s72[6]), .CP(clk), .CD(n1497), .Q(f72[6]) );
  CFD2QXL \f72_reg[5]  ( .D(s72[5]), .CP(clk), .CD(n1499), .Q(f72[5]) );
  CFD2QXL \f72_reg[2]  ( .D(s72[2]), .CP(clk), .CD(n1437), .Q(f72[2]) );
  CFD2QXL \f32_reg[9]  ( .D(w8[9]), .CP(clk), .CD(n1493), .Q(f32[9]) );
  CFD2QXL \f46_reg[9]  ( .D(n825), .CP(clk), .CD(n1453), .Q(f46[9]) );
  CFD2QXL \f53_reg[9]  ( .D(w11[9]), .CP(clk), .CD(n1462), .Q(f53[9]) );
  CFD2QXL \f63_reg[9]  ( .D(n827), .CP(clk), .CD(n1493), .Q(f63[9]) );
  CFD2QXL \f03_reg[31]  ( .D(n829), .CP(clk), .CD(n1464), .Q(f03[31]) );
  CFD2QXL \f36_reg[28]  ( .D(n830), .CP(clk), .CD(n1444), .Q(f36[28]) );
  CFD2QXL \f21_reg[15]  ( .D(n199), .CP(clk), .CD(n1431), .Q(f21[15]) );
  CFD2QXL \f21_reg[14]  ( .D(n821), .CP(clk), .CD(n1432), .Q(f21[14]) );
  CFD2QXL \f21_reg[13]  ( .D(n812), .CP(clk), .CD(n1432), .Q(f21[13]) );
  CFD2QXL \f11_reg[11]  ( .D(n813), .CP(clk), .CD(n1434), .Q(f11[11]) );
  CFD2QXL \f21_reg[12]  ( .D(n798), .CP(clk), .CD(n1433), .Q(f21[12]) );
  CFD2QXL \f21_reg[11]  ( .D(n802), .CP(clk), .CD(n1433), .Q(f21[11]) );
  CFD2QXL \f21_reg[8]  ( .D(n794), .CP(clk), .CD(n1457), .Q(f21[8]) );
  CFD2QXL \f21_reg[7]  ( .D(n795), .CP(clk), .CD(n1458), .Q(f21[7]) );
  CFD2QXL \f21_reg[29]  ( .D(n789), .CP(clk), .CD(n1443), .Q(f21[29]) );
  CFD2QXL \f21_reg[28]  ( .D(n791), .CP(clk), .CD(n1444), .Q(f21[28]) );
  CFD2QXL \f36_reg[26]  ( .D(n793), .CP(clk), .CD(n1445), .Q(f36[26]) );
  CFD2QXL \f11_reg[27]  ( .D(n787), .CP(clk), .CD(n1445), .Q(f11[27]) );
  CFD2QXL \f11_reg[26]  ( .D(n788), .CP(clk), .CD(n1445), .Q(f11[26]) );
  CFD2QXL \captA_reg[22]  ( .D(n172), .CP(clk), .CD(n1427), .Q(captA[22]) );
  CFD2QXL \captB_reg[22]  ( .D(n140), .CP(clk), .CD(n1472), .Q(captB[22]) );
  CFD2QXL \captA_reg[21]  ( .D(n171), .CP(clk), .CD(n1427), .Q(captA[21]) );
  CFD2QXL \captB_reg[21]  ( .D(n139), .CP(clk), .CD(n1474), .Q(captB[21]) );
  CFD2QXL \captC_reg[21]  ( .D(n107), .CP(clk), .CD(n1447), .Q(captC[21]) );
  CFD2QXL \f36_reg[24]  ( .D(n786), .CP(clk), .CD(n1425), .Q(f36[24]) );
  CFD2QXL \f13_reg[0]  ( .D(n783), .CP(clk), .CD(n1441), .Q(f13[0]) );
  CFD2QXL \f36_reg[17]  ( .D(f21[17]), .CP(clk), .CD(n1429), .Q(f36[17]) );
  CFD2QXL \f36_reg[23]  ( .D(f21[23]), .CP(clk), .CD(n1425), .Q(f36[23]) );
  CFD2QXL \f36_reg[22]  ( .D(f21[22]), .CP(clk), .CD(n1426), .Q(f36[22]) );
  CFD2QXL \f03_reg[30]  ( .D(n779), .CP(clk), .CD(n1464), .Q(f03[30]) );
  CFD2QXL \f13_reg[29]  ( .D(n780), .CP(clk), .CD(n1482), .Q(f13[29]) );
  CFD2QXL \f13_reg[28]  ( .D(n198), .CP(clk), .CD(n1484), .Q(f13[28]) );
  CFD2QXL \f14_reg[30]  ( .D(w2[30]), .CP(clk), .CD(n1483), .Q(f14[30]) );
  CFD2QXL \f14_reg[28]  ( .D(w2[28]), .CP(clk), .CD(n1486), .Q(f14[28]) );
  CFD2QXL \f14_reg[26]  ( .D(w2[26]), .CP(clk), .CD(n1490), .Q(f14[26]) );
  CFD2QXL \f14_reg[8]  ( .D(w2[8]), .CP(clk), .CD(n1497), .Q(f14[8]) );
  CFD2QXL \f14_reg[4]  ( .D(w2[4]), .CP(clk), .CD(n1437), .Q(f14[4]) );
  CFD2QXL \f14_reg[10]  ( .D(w2[10]), .CP(clk), .CD(n1494), .Q(f14[10]) );
  CFD2QXL \f14_reg[6]  ( .D(w2[6]), .CP(clk), .CD(n1500), .Q(f14[6]) );
  CFD2QXL \f36_reg[27]  ( .D(n778), .CP(clk), .CD(n1445), .Q(f36[27]) );
  CFD2QXL \f36_reg[19]  ( .D(f21[19]), .CP(clk), .CD(n1428), .Q(f36[19]) );
  CFD2QXL \f36_reg[18]  ( .D(f21[18]), .CP(clk), .CD(n1429), .Q(f36[18]) );
  CFD2QXL \f21_reg[27]  ( .D(n197), .CP(clk), .CD(n1445), .Q(f21[27]) );
  CFD2QXL \f21_reg[26]  ( .D(n777), .CP(clk), .CD(n1445), .Q(f21[26]) );
  CFD2QXL \f36_reg[25]  ( .D(f21[25]), .CP(clk), .CD(n1424), .Q(f36[25]) );
  CFD2QXL \f36_reg[16]  ( .D(f21[16]), .CP(clk), .CD(n1430), .Q(f36[16]) );
  CFD2QXL \f21_reg[24]  ( .D(n196), .CP(clk), .CD(n1425), .Q(f21[24]) );
  CFD2QXL \f21_reg[17]  ( .D(n774), .CP(clk), .CD(n1430), .Q(f21[17]) );
  CFD2QXL \f21_reg[20]  ( .D(n771), .CP(clk), .CD(n1427), .Q(f21[20]) );
  CFD2QXL \f21_reg[23]  ( .D(n195), .CP(clk), .CD(n1425), .Q(f21[23]) );
  CFD2QXL \f13_reg[27]  ( .D(n764), .CP(clk), .CD(n1485), .Q(f13[27]) );
  CFD2QXL \f13_reg[26]  ( .D(n765), .CP(clk), .CD(n1487), .Q(f13[26]) );
  CFD2QXL \f21_reg[19]  ( .D(n767), .CP(clk), .CD(n1428), .Q(f21[19]) );
  CFD2QXL \f14_reg[24]  ( .D(w2[24]), .CP(clk), .CD(n1471), .Q(f14[24]) );
  CFD2QXL \f14_reg[22]  ( .D(w2[22]), .CP(clk), .CD(n1474), .Q(f14[22]) );
  CFD2QXL \f14_reg[20]  ( .D(w2[20]), .CP(clk), .CD(n1477), .Q(f14[20]) );
  CFD2QXL \f14_reg[18]  ( .D(w2[18]), .CP(clk), .CD(n1502), .Q(f14[18]) );
  CFD2QXL \f14_reg[16]  ( .D(w2[16]), .CP(clk), .CD(n1505), .Q(f14[16]) );
  CFD2QXL \f11_reg[23]  ( .D(n761), .CP(clk), .CD(n1426), .Q(f11[23]) );
  CFD2QXL \f03_reg[29]  ( .D(n756), .CP(clk), .CD(n1465), .Q(f03[29]) );
  CFD2QXL \f03_reg[28]  ( .D(n758), .CP(clk), .CD(n1465), .Q(f03[28]) );
  CFD2QXL \f02_reg[30]  ( .D(n760), .CP(clk), .CD(n1481), .Q(f02[30]) );
  CFD2QXL \f21_reg[18]  ( .D(n754), .CP(clk), .CD(n1429), .Q(f21[18]) );
  CFD2QXL \f21_reg[25]  ( .D(n192), .CP(clk), .CD(n1424), .Q(f21[25]) );
  CFD2QXL \f21_reg[16]  ( .D(n749), .CP(clk), .CD(n1430), .Q(f21[16]) );
  CFD2QXL \f21_reg[22]  ( .D(n751), .CP(clk), .CD(n1426), .Q(f21[22]) );
  CFD2QXL \f36_reg[21]  ( .D(f21[21]), .CP(clk), .CD(n1427), .Q(f36[21]) );
  CFD2QXL \f36_reg[20]  ( .D(f21[20]), .CP(clk), .CD(n1427), .Q(f36[20]) );
  CFD2QXL \f14_reg[31]  ( .D(w2[31]), .CP(clk), .CD(n1481), .Q(f14[31]) );
  CFD2QXL \f13_reg[25]  ( .D(n743), .CP(clk), .CD(n1489), .Q(f13[25]) );
  CFD2QXL \f13_reg[24]  ( .D(n745), .CP(clk), .CD(n1468), .Q(f13[24]) );
  CFD2QXL \f21_reg[21]  ( .D(n747), .CP(clk), .CD(n1427), .Q(f21[21]) );
  CFD2QXL \f12_reg[30]  ( .D(w1[30]), .CP(clk), .CD(n1444), .Q(f12[30]) );
  CFD2QXL \f01_reg[30]  ( .D(n738), .CP(clk), .CD(n1443), .Q(f01[30]) );
  CFD2QXL \f01_reg[28]  ( .D(n739), .CP(clk), .CD(n1444), .Q(f01[28]) );
  CFD2QXL \f01_reg[26]  ( .D(n741), .CP(clk), .CD(n1424), .Q(f01[26]) );
  CFD2QXL \f01_reg[24]  ( .D(n729), .CP(clk), .CD(n1425), .Q(f01[24]) );
  CFD2QXL \f01_reg[22]  ( .D(n731), .CP(clk), .CD(n1426), .Q(f01[22]) );
  CFD2QXL \f01_reg[18]  ( .D(n733), .CP(clk), .CD(n1429), .Q(f01[18]) );
  CFD2QXL \f03_reg[26]  ( .D(n727), .CP(clk), .CD(n1466), .Q(f03[26]) );
  CFD2QXL \f02_reg[31]  ( .D(n724), .CP(clk), .CD(n1480), .Q(f02[31]) );
  CFD2QXL \f13_reg[22]  ( .D(n725), .CP(clk), .CD(n1471), .Q(f13[22]) );
  CFD2QXL \f03_reg[27]  ( .D(n722), .CP(clk), .CD(n1466), .Q(f03[27]) );
  CFD2QXL \f12_reg[31]  ( .D(w1[31]), .CP(clk), .CD(n1443), .Q(f12[31]) );
  CFD2QXL \f13_reg[20]  ( .D(n718), .CP(clk), .CD(n1474), .Q(f13[20]) );
  CFD2QX1 \f03_reg[10]  ( .D(n720), .CP(clk), .CD(n1452), .Q(f03[10]) );
  CFD2QXL \f14_reg[29]  ( .D(w2[29]), .CP(clk), .CD(n1485), .Q(f14[29]) );
  CFD2QXL \f01_reg[31]  ( .D(n717), .CP(clk), .CD(n1442), .Q(f01[31]) );
  CFD2QXL \f13_reg[18]  ( .D(n713), .CP(clk), .CD(n1511), .Q(f13[18]) );
  CFD2QXL \f13_reg[16]  ( .D(n715), .CP(clk), .CD(n1511), .Q(f13[16]) );
  CFD2QXL \f15_reg[31]  ( .D(w3[31]), .CP(clk), .CD(n1465), .Q(f15[31]) );
  CFD2QXL \f15_reg[23]  ( .D(w3[23]), .CP(clk), .CD(n1446), .Q(f15[23]) );
  CFD2QXL \f15_reg[22]  ( .D(w3[22]), .CP(clk), .CD(n1447), .Q(f15[22]) );
  CFD2QXL \f15_reg[21]  ( .D(w3[21]), .CP(clk), .CD(n1447), .Q(f15[21]) );
  CFD2QXL \f15_reg[20]  ( .D(w3[20]), .CP(clk), .CD(n1448), .Q(f15[20]) );
  CFD2QXL \f15_reg[19]  ( .D(w3[19]), .CP(clk), .CD(n1448), .Q(f15[19]) );
  CFD2QXL \f15_reg[18]  ( .D(w3[18]), .CP(clk), .CD(n1449), .Q(f15[18]) );
  CFD2QXL \f15_reg[17]  ( .D(w3[17]), .CP(clk), .CD(n1449), .Q(f15[17]) );
  CFD2QXL \f15_reg[16]  ( .D(w3[16]), .CP(clk), .CD(n1450), .Q(f15[16]) );
  CFD2QXL \f15_reg[15]  ( .D(w3[15]), .CP(clk), .CD(n1450), .Q(f15[15]) );
  CFD2QXL \f15_reg[14]  ( .D(w3[14]), .CP(clk), .CD(n1450), .Q(f15[14]) );
  CFD2QXL \f15_reg[13]  ( .D(w3[13]), .CP(clk), .CD(n1451), .Q(f15[13]) );
  CFD2QXL \f15_reg[12]  ( .D(w3[12]), .CP(clk), .CD(n1451), .Q(f15[12]) );
  CFD2QXL \f15_reg[11]  ( .D(w3[11]), .CP(clk), .CD(n1452), .Q(f15[11]) );
  CFD2QXL \f26_reg[9]  ( .D(w4[9]), .CP(clk), .CD(n1457), .Q(f26[9]) );
  CFD2QXL \f26_reg[8]  ( .D(w4[8]), .CP(clk), .CD(n1458), .Q(f26[8]) );
  CFD2QXL \f26_reg[7]  ( .D(w4[7]), .CP(clk), .CD(n1458), .Q(f26[7]) );
  CFD2QXL \f28_reg[8]  ( .D(w6[8]), .CP(clk), .CD(n1495), .Q(f28[8]) );
  CFD2QXL \f28_reg[7]  ( .D(w6[7]), .CP(clk), .CD(n1496), .Q(f28[7]) );
  CFD2QXL \f28_reg[6]  ( .D(w6[6]), .CP(clk), .CD(n1498), .Q(f28[6]) );
  CFD2QXL \f31_reg[5]  ( .D(w7[5]), .CP(clk), .CD(n1500), .Q(f31[5]) );
  CFD2QXL \f31_reg[4]  ( .D(w7[4]), .CP(clk), .CD(n1435), .Q(f31[4]) );
  CFD2QXL \f31_reg[3]  ( .D(w7[3]), .CP(clk), .CD(n1437), .Q(f31[3]) );
  CFD2QXL \f41_reg[31]  ( .D(s41[31]), .CP(clk), .CD(n1479), .Q(f41[31]) );
  CFD2QXL \f41_reg[30]  ( .D(s41[30]), .CP(clk), .CD(n1481), .Q(f41[30]) );
  CFD2QXL \f41_reg[0]  ( .D(s41[0]), .CP(clk), .CD(n1441), .Q(f41[0]) );
  CFD2QXL \f42_reg[31]  ( .D(s42[31]), .CP(clk), .CD(n1479), .Q(f42[31]) );
  CFD2QXL \f42_reg[30]  ( .D(s42[30]), .CP(clk), .CD(n1480), .Q(f42[30]) );
  CFD2QXL \f42_reg[0]  ( .D(s42[0]), .CP(clk), .CD(n1440), .Q(f42[0]) );
  CFD2QXL \f54_reg[31]  ( .D(s54[31]), .CP(clk), .CD(n1480), .Q(f54[31]) );
  CFD2QXL \f54_reg[30]  ( .D(s54[30]), .CP(clk), .CD(n1481), .Q(f54[30]) );
  CFD2QXL \f54_reg[1]  ( .D(s54[1]), .CP(clk), .CD(n1440), .Q(f54[1]) );
  CFD2QXL \f54_reg[0]  ( .D(s54[0]), .CP(clk), .CD(n1441), .Q(f54[0]) );
  CFD2QXL \f61_reg[31]  ( .D(s61[31]), .CP(clk), .CD(n1479), .Q(f61[31]) );
  CFD2QXL \f61_reg[30]  ( .D(s61[30]), .CP(clk), .CD(n1481), .Q(f61[30]) );
  CFD2QXL \f61_reg[0]  ( .D(s61[0]), .CP(clk), .CD(n1441), .Q(f61[0]) );
  CFD2QXL all_in_reg ( .D(N7), .CP(clk), .CD(n1464), .Q(all_in) );
  CFD2QXL all_in1_reg ( .D(n269), .CP(clk), .CD(n1464), .Q(all_in1) );
  CFD2QXL all_in2_reg ( .D(n267), .CP(clk), .CD(n1464), .Q(all_in2) );
  CFD2QXL all_in3_reg ( .D(n642), .CP(clk), .CD(n1464), .Q(all_in3) );
  CFD2QXL all_in4_reg ( .D(n644), .CP(clk), .CD(n1464), .Q(all_in4) );
  CFD2QXL all_in5_reg ( .D(n646), .CP(clk), .CD(n1464), .Q(all_in5) );
  CFD2QXL all_in6_reg ( .D(n285), .CP(clk), .CD(n1464), .Q(all_in6) );
  CFD2QXL all_in7_reg ( .D(n648), .CP(clk), .CD(n1464), .Q(all_in7) );
  CFD2QXL all_in8_reg ( .D(n638), .CP(clk), .CD(n1463), .Q(all_in8) );
  CFD2QXL all_in9_reg ( .D(n640), .CP(clk), .CD(n1463), .Q(all_in9) );
  CFD2QXL \f15_reg[30]  ( .D(w3[30]), .CP(clk), .CD(n1465), .Q(f15[30]) );
  CFD2QXL \f15_reg[29]  ( .D(w3[29]), .CP(clk), .CD(n1466), .Q(f15[29]) );
  CFD2QXL \f15_reg[28]  ( .D(w3[28]), .CP(clk), .CD(n1466), .Q(f15[28]) );
  CFD2QXL \f15_reg[27]  ( .D(w3[27]), .CP(clk), .CD(n1466), .Q(f15[27]) );
  CFD2QXL \f15_reg[26]  ( .D(w3[26]), .CP(clk), .CD(n1467), .Q(f15[26]) );
  CFD2QXL \f15_reg[25]  ( .D(w3[25]), .CP(clk), .CD(n1467), .Q(f15[25]) );
  CFD2QXL \f15_reg[24]  ( .D(w3[24]), .CP(clk), .CD(n1446), .Q(f15[24]) );
  CFD2QXL \f15_reg[10]  ( .D(w3[10]), .CP(clk), .CD(n1452), .Q(f15[10]) );
  CFD2QXL \f15_reg[9]  ( .D(w3[9]), .CP(clk), .CD(n1453), .Q(f15[9]) );
  CFD2QXL \f15_reg[8]  ( .D(w3[8]), .CP(clk), .CD(n1453), .Q(f15[8]) );
  CFD2QXL \f15_reg[7]  ( .D(w3[7]), .CP(clk), .CD(n1454), .Q(f15[7]) );
  CFD2QXL \f15_reg[6]  ( .D(w3[6]), .CP(clk), .CD(n1454), .Q(f15[6]) );
  CFD2QXL \f15_reg[5]  ( .D(w3[5]), .CP(clk), .CD(n1455), .Q(f15[5]) );
  CFD2QXL \f15_reg[4]  ( .D(w3[4]), .CP(clk), .CD(n1455), .Q(f15[4]) );
  CFD2QXL \f15_reg[3]  ( .D(w3[3]), .CP(clk), .CD(n1456), .Q(f15[3]) );
  CFD2QXL \f15_reg[2]  ( .D(w3[2]), .CP(clk), .CD(n1456), .Q(f15[2]) );
  CFD2QXL \f15_reg[0]  ( .D(w3[0]), .CP(clk), .CD(n1456), .Q(f15[0]) );
  CFD2QXL \f23_reg[31]  ( .D(n636), .CP(clk), .CD(n1465), .Q(f23[31]) );
  CFD2QXL \f23_reg[30]  ( .D(n628), .CP(clk), .CD(n1465), .Q(f23[30]) );
  CFD2QXL \f23_reg[29]  ( .D(n630), .CP(clk), .CD(n1465), .Q(f23[29]) );
  CFD2QXL \f23_reg[28]  ( .D(n632), .CP(clk), .CD(n1466), .Q(f23[28]) );
  CFD2QXL \f23_reg[27]  ( .D(n287), .CP(clk), .CD(n1466), .Q(f23[27]) );
  CFD2QXL \f23_reg[26]  ( .D(n634), .CP(clk), .CD(n1467), .Q(f23[26]) );
  CFD2QXL \f23_reg[25]  ( .D(n620), .CP(clk), .CD(n1467), .Q(f23[25]) );
  CFD2QXL \f23_reg[24]  ( .D(n622), .CP(clk), .CD(n1446), .Q(f23[24]) );
  CFD2QXL \f23_reg[23]  ( .D(n624), .CP(clk), .CD(n1446), .Q(f23[23]) );
  CFD2QXL \f23_reg[22]  ( .D(n289), .CP(clk), .CD(n1447), .Q(f23[22]) );
  CFD2QXL \f23_reg[21]  ( .D(n626), .CP(clk), .CD(n1447), .Q(f23[21]) );
  CFD2QXL \f23_reg[20]  ( .D(n612), .CP(clk), .CD(n1448), .Q(f23[20]) );
  CFD2QXL \f23_reg[19]  ( .D(n614), .CP(clk), .CD(n1448), .Q(f23[19]) );
  CFD2QXL \f23_reg[18]  ( .D(n616), .CP(clk), .CD(n1449), .Q(f23[18]) );
  CFD2QXL \f23_reg[17]  ( .D(n291), .CP(clk), .CD(n1449), .Q(f23[17]) );
  CFD2QXL \f23_reg[16]  ( .D(n618), .CP(clk), .CD(n1449), .Q(f23[16]) );
  CFD2QXL \f23_reg[15]  ( .D(n604), .CP(clk), .CD(n1450), .Q(f23[15]) );
  CFD2QXL \f23_reg[14]  ( .D(n606), .CP(clk), .CD(n1450), .Q(f23[14]) );
  CFD2QXL \f23_reg[13]  ( .D(n608), .CP(clk), .CD(n1451), .Q(f23[13]) );
  CFD2QXL \f23_reg[12]  ( .D(n293), .CP(clk), .CD(n1451), .Q(f23[12]) );
  CFD2QXL \f23_reg[11]  ( .D(n610), .CP(clk), .CD(n1452), .Q(f23[11]) );
  CFD2QXL \f23_reg[10]  ( .D(n596), .CP(clk), .CD(n1452), .Q(f23[10]) );
  CFD2QXL \f23_reg[9]  ( .D(n598), .CP(clk), .CD(n1453), .Q(f23[9]) );
  CFD2QXL \f23_reg[8]  ( .D(n600), .CP(clk), .CD(n1453), .Q(f23[8]) );
  CFD2QXL \f23_reg[7]  ( .D(n295), .CP(clk), .CD(n1454), .Q(f23[7]) );
  CFD2QXL \f23_reg[6]  ( .D(n602), .CP(clk), .CD(n1454), .Q(f23[6]) );
  CFD2QXL \f23_reg[5]  ( .D(n588), .CP(clk), .CD(n1455), .Q(f23[5]) );
  CFD2QXL \f23_reg[4]  ( .D(n590), .CP(clk), .CD(n1455), .Q(f23[4]) );
  CFD2QXL \f23_reg[3]  ( .D(n592), .CP(clk), .CD(n1455), .Q(f23[3]) );
  CFD2QXL \f23_reg[2]  ( .D(n297), .CP(clk), .CD(n1456), .Q(f23[2]) );
  CFD2QXL \f23_reg[0]  ( .D(n594), .CP(clk), .CD(n1456), .Q(f23[0]) );
  CFD2QXL \f26_reg[31]  ( .D(w4[31]), .CP(clk), .CD(n1442), .Q(f26[31]) );
  CFD2QXL \f26_reg[30]  ( .D(w4[30]), .CP(clk), .CD(n1443), .Q(f26[30]) );
  CFD2QXL \f26_reg[29]  ( .D(w4[29]), .CP(clk), .CD(n1443), .Q(f26[29]) );
  CFD2QXL \f26_reg[28]  ( .D(w4[28]), .CP(clk), .CD(n1444), .Q(f26[28]) );
  CFD2QXL \f26_reg[27]  ( .D(w4[27]), .CP(clk), .CD(n1445), .Q(f26[27]) );
  CFD2QXL \f26_reg[26]  ( .D(w4[26]), .CP(clk), .CD(n1429), .Q(f26[26]) );
  CFD2QXL \f26_reg[25]  ( .D(w4[25]), .CP(clk), .CD(n1424), .Q(f26[25]) );
  CFD2QXL \f26_reg[24]  ( .D(w4[24]), .CP(clk), .CD(n1425), .Q(f26[24]) );
  CFD2QXL \f26_reg[23]  ( .D(w4[23]), .CP(clk), .CD(n1426), .Q(f26[23]) );
  CFD2QXL \f26_reg[22]  ( .D(w4[22]), .CP(clk), .CD(n1426), .Q(f26[22]) );
  CFD2QXL \f26_reg[21]  ( .D(w4[21]), .CP(clk), .CD(n1427), .Q(f26[21]) );
  CFD2QXL \f26_reg[20]  ( .D(w4[20]), .CP(clk), .CD(n1428), .Q(f26[20]) );
  CFD2QXL \f26_reg[19]  ( .D(w4[19]), .CP(clk), .CD(n1428), .Q(f26[19]) );
  CFD2QXL \f26_reg[18]  ( .D(w4[18]), .CP(clk), .CD(n1429), .Q(f26[18]) );
  CFD2QXL \f26_reg[17]  ( .D(w4[17]), .CP(clk), .CD(n1430), .Q(f26[17]) );
  CFD2QXL \f26_reg[16]  ( .D(w4[16]), .CP(clk), .CD(n1430), .Q(f26[16]) );
  CFD2QXL \f26_reg[15]  ( .D(w4[15]), .CP(clk), .CD(n1431), .Q(f26[15]) );
  CFD2QXL \f26_reg[14]  ( .D(w4[14]), .CP(clk), .CD(n1432), .Q(f26[14]) );
  CFD2QXL \f26_reg[13]  ( .D(w4[13]), .CP(clk), .CD(n1432), .Q(f26[13]) );
  CFD2QXL \f26_reg[12]  ( .D(w4[12]), .CP(clk), .CD(n1433), .Q(f26[12]) );
  CFD2QXL \f26_reg[11]  ( .D(w4[11]), .CP(clk), .CD(n1434), .Q(f26[11]) );
  CFD2QXL \f26_reg[10]  ( .D(w4[10]), .CP(clk), .CD(n1434), .Q(f26[10]) );
  CFD2QXL \f26_reg[6]  ( .D(w4[6]), .CP(clk), .CD(n1459), .Q(f26[6]) );
  CFD2QXL \f26_reg[5]  ( .D(w4[5]), .CP(clk), .CD(n1460), .Q(f26[5]) );
  CFD2QXL \f26_reg[4]  ( .D(w4[4]), .CP(clk), .CD(n1460), .Q(f26[4]) );
  CFD2QXL \f26_reg[3]  ( .D(w4[3]), .CP(clk), .CD(n1461), .Q(f26[3]) );
  CFD2QXL \f26_reg[2]  ( .D(w4[2]), .CP(clk), .CD(n1462), .Q(f26[2]) );
  CFD2QXL \f26_reg[1]  ( .D(w4[1]), .CP(clk), .CD(n1462), .Q(f26[1]) );
  CFD2QXL \f26_reg[0]  ( .D(w4[0]), .CP(clk), .CD(n1463), .Q(f26[0]) );
  CFD2QXL \f28_reg[31]  ( .D(w6[31]), .CP(clk), .CD(n1479), .Q(f28[31]) );
  CFD2QXL \f28_reg[30]  ( .D(w6[30]), .CP(clk), .CD(n1481), .Q(f28[30]) );
  CFD2QXL \f28_reg[29]  ( .D(w6[29]), .CP(clk), .CD(n1482), .Q(f28[29]) );
  CFD2QXL \f28_reg[28]  ( .D(w6[28]), .CP(clk), .CD(n1484), .Q(f28[28]) );
  CFD2QXL \f28_reg[27]  ( .D(w6[27]), .CP(clk), .CD(n1486), .Q(f28[27]) );
  CFD2QXL \f28_reg[26]  ( .D(w6[26]), .CP(clk), .CD(n1487), .Q(f28[26]) );
  CFD2QXL \f28_reg[25]  ( .D(w6[25]), .CP(clk), .CD(n1489), .Q(f28[25]) );
  CFD2QXL \f28_reg[24]  ( .D(w6[24]), .CP(clk), .CD(n1468), .Q(f28[24]) );
  CFD2QXL \f28_reg[23]  ( .D(w6[23]), .CP(clk), .CD(n1470), .Q(f28[23]) );
  CFD2QXL \f28_reg[22]  ( .D(w6[22]), .CP(clk), .CD(n1471), .Q(f28[22]) );
  CFD2QXL \f28_reg[21]  ( .D(w6[21]), .CP(clk), .CD(n1473), .Q(f28[21]) );
  CFD2QXL \f28_reg[20]  ( .D(w6[20]), .CP(clk), .CD(n1475), .Q(f28[20]) );
  CFD2QXL \f28_reg[19]  ( .D(w6[19]), .CP(clk), .CD(n1476), .Q(f28[19]) );
  CFD2QXL \f28_reg[18]  ( .D(w6[18]), .CP(clk), .CD(n1478), .Q(f28[18]) );
  CFD2QXL \f28_reg[17]  ( .D(w6[17]), .CP(clk), .CD(n1501), .Q(f28[17]) );
  CFD2QXL \f28_reg[16]  ( .D(w6[16]), .CP(clk), .CD(n1503), .Q(f28[16]) );
  CFD2QXL \f28_reg[15]  ( .D(w6[15]), .CP(clk), .CD(n1504), .Q(f28[15]) );
  CFD2QXL \f28_reg[14]  ( .D(w6[14]), .CP(clk), .CD(n1506), .Q(f28[14]) );
  CFD2QXL \f28_reg[13]  ( .D(w6[13]), .CP(clk), .CD(n1507), .Q(f28[13]) );
  CFD2QXL \f28_reg[12]  ( .D(w6[12]), .CP(clk), .CD(n1509), .Q(f28[12]) );
  CFD2QXL \f28_reg[11]  ( .D(w6[11]), .CP(clk), .CD(n1490), .Q(f28[11]) );
  CFD2QXL \f28_reg[10]  ( .D(w6[10]), .CP(clk), .CD(n1491), .Q(f28[10]) );
  CFD2QXL \f28_reg[9]  ( .D(w6[9]), .CP(clk), .CD(n1493), .Q(f28[9]) );
  CFD2QXL \f28_reg[5]  ( .D(w6[5]), .CP(clk), .CD(n1499), .Q(f28[5]) );
  CFD2QXL \f28_reg[4]  ( .D(w6[4]), .CP(clk), .CD(n1435), .Q(f28[4]) );
  CFD2QXL \f28_reg[3]  ( .D(w6[3]), .CP(clk), .CD(n1436), .Q(f28[3]) );
  CFD2QXL \f28_reg[2]  ( .D(w6[2]), .CP(clk), .CD(n1438), .Q(f28[2]) );
  CFD2QXL \f28_reg[1]  ( .D(w6[1]), .CP(clk), .CD(n1439), .Q(f28[1]) );
  CFD2QXL \f28_reg[0]  ( .D(w6[0]), .CP(clk), .CD(n1441), .Q(f28[0]) );
  CFD2QXL \f31_reg[31]  ( .D(w7[31]), .CP(clk), .CD(n1480), .Q(f31[31]) );
  CFD2QXL \f31_reg[29]  ( .D(w7[29]), .CP(clk), .CD(n1483), .Q(f31[29]) );
  CFD2QXL \f31_reg[28]  ( .D(w7[28]), .CP(clk), .CD(n1485), .Q(f31[28]) );
  CFD2QXL \f31_reg[27]  ( .D(w7[27]), .CP(clk), .CD(n1486), .Q(f31[27]) );
  CFD2QXL \f31_reg[26]  ( .D(w7[26]), .CP(clk), .CD(n1488), .Q(f31[26]) );
  CFD2QXL \f31_reg[25]  ( .D(w7[25]), .CP(clk), .CD(n1489), .Q(f31[25]) );
  CFD2QXL \f31_reg[24]  ( .D(w7[24]), .CP(clk), .CD(n1469), .Q(f31[24]) );
  CFD2QXL \f31_reg[23]  ( .D(w7[23]), .CP(clk), .CD(n1470), .Q(f31[23]) );
  CFD2QXL \f31_reg[22]  ( .D(w7[22]), .CP(clk), .CD(n1472), .Q(f31[22]) );
  CFD2QXL \f31_reg[21]  ( .D(w7[21]), .CP(clk), .CD(n1474), .Q(f31[21]) );
  CFD2QXL \f31_reg[20]  ( .D(w7[20]), .CP(clk), .CD(n1475), .Q(f31[20]) );
  CFD2QXL \f31_reg[19]  ( .D(w7[19]), .CP(clk), .CD(n1477), .Q(f31[19]) );
  CFD2QXL \f31_reg[18]  ( .D(w7[18]), .CP(clk), .CD(n1478), .Q(f31[18]) );
  CFD2QXL \f31_reg[17]  ( .D(w7[17]), .CP(clk), .CD(n1502), .Q(f31[17]) );
  CFD2QXL \f31_reg[16]  ( .D(w7[16]), .CP(clk), .CD(n1503), .Q(f31[16]) );
  CFD2QXL \f31_reg[15]  ( .D(w7[15]), .CP(clk), .CD(n1505), .Q(f31[15]) );
  CFD2QXL \f31_reg[14]  ( .D(w7[14]), .CP(clk), .CD(n1506), .Q(f31[14]) );
  CFD2QXL \f31_reg[13]  ( .D(w7[13]), .CP(clk), .CD(n1508), .Q(f31[13]) );
  CFD2QXL \f31_reg[12]  ( .D(w7[12]), .CP(clk), .CD(n1509), .Q(f31[12]) );
  CFD2QXL \f31_reg[11]  ( .D(w7[11]), .CP(clk), .CD(n1491), .Q(f31[11]) );
  CFD2QXL \f31_reg[10]  ( .D(w7[10]), .CP(clk), .CD(n1492), .Q(f31[10]) );
  CFD2QXL \f31_reg[9]  ( .D(w7[9]), .CP(clk), .CD(n1494), .Q(f31[9]) );
  CFD2QXL \f31_reg[8]  ( .D(w7[8]), .CP(clk), .CD(n1495), .Q(f31[8]) );
  CFD2QXL \f31_reg[7]  ( .D(w7[7]), .CP(clk), .CD(n1497), .Q(f31[7]) );
  CFD2QXL \f31_reg[6]  ( .D(w7[6]), .CP(clk), .CD(n1499), .Q(f31[6]) );
  CFD2QXL \f31_reg[2]  ( .D(w7[2]), .CP(clk), .CD(n1438), .Q(f31[2]) );
  CFD2QXL \f31_reg[1]  ( .D(w7[1]), .CP(clk), .CD(n1440), .Q(f31[1]) );
  CFD2QXL \f31_reg[0]  ( .D(w7[0]), .CP(clk), .CD(n1441), .Q(f31[0]) );
  CFD2QXL \f37_reg[31]  ( .D(n584), .CP(clk), .CD(n1464), .Q(f37[31]) );
  CFD2QXL \f37_reg[30]  ( .D(n299), .CP(clk), .CD(n1465), .Q(f37[30]) );
  CFD2QXL \f37_reg[29]  ( .D(n586), .CP(clk), .CD(n1465), .Q(f37[29]) );
  CFD2QXL \f37_reg[28]  ( .D(n576), .CP(clk), .CD(n1466), .Q(f37[28]) );
  CFD2QXL \f37_reg[27]  ( .D(n578), .CP(clk), .CD(n1466), .Q(f37[27]) );
  CFD2QXL \f37_reg[26]  ( .D(n580), .CP(clk), .CD(n1467), .Q(f37[26]) );
  CFD2QXL \f37_reg[25]  ( .D(n301), .CP(clk), .CD(n1467), .Q(f37[25]) );
  CFD2QXL \f37_reg[24]  ( .D(n582), .CP(clk), .CD(n1446), .Q(f37[24]) );
  CFD2QXL \f37_reg[23]  ( .D(n568), .CP(clk), .CD(n1446), .Q(f37[23]) );
  CFD2QXL \f37_reg[22]  ( .D(n570), .CP(clk), .CD(n1447), .Q(f37[22]) );
  CFD2QXL \f37_reg[21]  ( .D(n572), .CP(clk), .CD(n1447), .Q(f37[21]) );
  CFD2QXL \f37_reg[20]  ( .D(n303), .CP(clk), .CD(n1448), .Q(f37[20]) );
  CFD2QXL \f37_reg[19]  ( .D(n574), .CP(clk), .CD(n1448), .Q(f37[19]) );
  CFD2QXL \f37_reg[18]  ( .D(n434), .CP(clk), .CD(n1448), .Q(f37[18]) );
  CFD2QXL \f37_reg[17]  ( .D(n436), .CP(clk), .CD(n1449), .Q(f37[17]) );
  CFD2QXL \f37_reg[16]  ( .D(n336), .CP(clk), .CD(n1449), .Q(f37[16]) );
  CFD2QXL \f37_reg[15]  ( .D(n305), .CP(clk), .CD(n1450), .Q(f37[15]) );
  CFD2QXL \f37_reg[14]  ( .D(n566), .CP(clk), .CD(n1450), .Q(f37[14]) );
  CFD2QXL \f37_reg[13]  ( .D(n426), .CP(clk), .CD(n1451), .Q(f37[13]) );
  CFD2QXL \f37_reg[12]  ( .D(n428), .CP(clk), .CD(n1451), .Q(f37[12]) );
  CFD2QXL \f37_reg[11]  ( .D(n338), .CP(clk), .CD(n1452), .Q(f37[11]) );
  CFD2QXL \f37_reg[10]  ( .D(n430), .CP(clk), .CD(n1452), .Q(f37[10]) );
  CFD2QXL \f37_reg[9]  ( .D(n432), .CP(clk), .CD(n1453), .Q(f37[9]) );
  CFD2QXL \f37_reg[8]  ( .D(n418), .CP(clk), .CD(n1453), .Q(f37[8]) );
  CFD2QXL \f37_reg[7]  ( .D(n420), .CP(clk), .CD(n1454), .Q(f37[7]) );
  CFD2QXL \f37_reg[6]  ( .D(n340), .CP(clk), .CD(n1454), .Q(f37[6]) );
  CFD2QXL \f37_reg[5]  ( .D(n422), .CP(clk), .CD(n1454), .Q(f37[5]) );
  CFD2QXL \f37_reg[4]  ( .D(n424), .CP(clk), .CD(n1455), .Q(f37[4]) );
  CFD2QXL \f37_reg[3]  ( .D(n414), .CP(clk), .CD(n1455), .Q(f37[3]) );
  CFD2QXL \f37_reg[2]  ( .D(n416), .CP(clk), .CD(n1456), .Q(f37[2]) );
  CFD2QXL \f37_reg[0]  ( .D(n342), .CP(clk), .CD(n1456), .Q(f37[0]) );
  CFD2QXL \f41_reg[29]  ( .D(s41[29]), .CP(clk), .CD(n1483), .Q(f41[29]) );
  CFD2QXL \f41_reg[28]  ( .D(s41[28]), .CP(clk), .CD(n1484), .Q(f41[28]) );
  CFD2QXL \f41_reg[27]  ( .D(s41[27]), .CP(clk), .CD(n1486), .Q(f41[27]) );
  CFD2QXL \f41_reg[26]  ( .D(s41[26]), .CP(clk), .CD(n1487), .Q(f41[26]) );
  CFD2QXL \f41_reg[25]  ( .D(s41[25]), .CP(clk), .CD(n1489), .Q(f41[25]) );
  CFD2QXL \f41_reg[24]  ( .D(s41[24]), .CP(clk), .CD(n1468), .Q(f41[24]) );
  CFD2QXL \f41_reg[23]  ( .D(s41[23]), .CP(clk), .CD(n1470), .Q(f41[23]) );
  CFD2QXL \f41_reg[22]  ( .D(s41[22]), .CP(clk), .CD(n1472), .Q(f41[22]) );
  CFD2QXL \f41_reg[21]  ( .D(s41[21]), .CP(clk), .CD(n1473), .Q(f41[21]) );
  CFD2QXL \f41_reg[20]  ( .D(s41[20]), .CP(clk), .CD(n1475), .Q(f41[20]) );
  CFD2QXL \f41_reg[19]  ( .D(s41[19]), .CP(clk), .CD(n1476), .Q(f41[19]) );
  CFD2QXL \f41_reg[18]  ( .D(s41[18]), .CP(clk), .CD(n1478), .Q(f41[18]) );
  CFD2QXL \f41_reg[17]  ( .D(s41[17]), .CP(clk), .CD(n1502), .Q(f41[17]) );
  CFD2QXL \f41_reg[16]  ( .D(s41[16]), .CP(clk), .CD(n1503), .Q(f41[16]) );
  CFD2QXL \f41_reg[15]  ( .D(s41[15]), .CP(clk), .CD(n1505), .Q(f41[15]) );
  CFD2QXL \f41_reg[14]  ( .D(s41[14]), .CP(clk), .CD(n1506), .Q(f41[14]) );
  CFD2QXL \f41_reg[13]  ( .D(s41[13]), .CP(clk), .CD(n1508), .Q(f41[13]) );
  CFD2QXL \f41_reg[12]  ( .D(s41[12]), .CP(clk), .CD(n1510), .Q(f41[12]) );
  CFD2QXL \f41_reg[11]  ( .D(s41[11]), .CP(clk), .CD(n1490), .Q(f41[11]) );
  CFD2QXL \f41_reg[10]  ( .D(s41[10]), .CP(clk), .CD(n1492), .Q(f41[10]) );
  CFD2QXL \f41_reg[9]  ( .D(s41[9]), .CP(clk), .CD(n1493), .Q(f41[9]) );
  CFD2QXL \f41_reg[8]  ( .D(s41[8]), .CP(clk), .CD(n1495), .Q(f41[8]) );
  CFD2QXL \f41_reg[7]  ( .D(s41[7]), .CP(clk), .CD(n1497), .Q(f41[7]) );
  CFD2QXL \f41_reg[6]  ( .D(s41[6]), .CP(clk), .CD(n1498), .Q(f41[6]) );
  CFD2QXL \f41_reg[5]  ( .D(s41[5]), .CP(clk), .CD(n1500), .Q(f41[5]) );
  CFD2QXL \f41_reg[4]  ( .D(s41[4]), .CP(clk), .CD(n1435), .Q(f41[4]) );
  CFD2QXL \f41_reg[3]  ( .D(s41[3]), .CP(clk), .CD(n1436), .Q(f41[3]) );
  CFD2QXL \f41_reg[2]  ( .D(s41[2]), .CP(clk), .CD(n1438), .Q(f41[2]) );
  CFD2QXL \f41_reg[1]  ( .D(s41[1]), .CP(clk), .CD(n1439), .Q(f41[1]) );
  CFD2QXL \f42_reg[29]  ( .D(s42[29]), .CP(clk), .CD(n1482), .Q(f42[29]) );
  CFD2QXL \f42_reg[28]  ( .D(s42[28]), .CP(clk), .CD(n1484), .Q(f42[28]) );
  CFD2QXL \f42_reg[27]  ( .D(s42[27]), .CP(clk), .CD(n1485), .Q(f42[27]) );
  CFD2QXL \f42_reg[26]  ( .D(s42[26]), .CP(clk), .CD(n1487), .Q(f42[26]) );
  CFD2QXL \f42_reg[25]  ( .D(s42[25]), .CP(clk), .CD(n1488), .Q(f42[25]) );
  CFD2QXL \f42_reg[24]  ( .D(s42[24]), .CP(clk), .CD(n1468), .Q(f42[24]) );
  CFD2QXL \f42_reg[23]  ( .D(s42[23]), .CP(clk), .CD(n1469), .Q(f42[23]) );
  CFD2QXL \f42_reg[22]  ( .D(s42[22]), .CP(clk), .CD(n1471), .Q(f42[22]) );
  CFD2QXL \f42_reg[21]  ( .D(s42[21]), .CP(clk), .CD(n1473), .Q(f42[21]) );
  CFD2QXL \f42_reg[20]  ( .D(s42[20]), .CP(clk), .CD(n1474), .Q(f42[20]) );
  CFD2QXL \f42_reg[19]  ( .D(s42[19]), .CP(clk), .CD(n1476), .Q(f42[19]) );
  CFD2QXL \f42_reg[18]  ( .D(s42[18]), .CP(clk), .CD(n1477), .Q(f42[18]) );
  CFD2QXL \f42_reg[17]  ( .D(s42[17]), .CP(clk), .CD(n1501), .Q(f42[17]) );
  CFD2QXL \f42_reg[16]  ( .D(s42[16]), .CP(clk), .CD(n1503), .Q(f42[16]) );
  CFD2QXL \f42_reg[15]  ( .D(s42[15]), .CP(clk), .CD(n1504), .Q(f42[15]) );
  CFD2QXL \f42_reg[14]  ( .D(s42[14]), .CP(clk), .CD(n1506), .Q(f42[14]) );
  CFD2QXL \f42_reg[13]  ( .D(s42[13]), .CP(clk), .CD(n1507), .Q(f42[13]) );
  CFD2QXL \f42_reg[12]  ( .D(s42[12]), .CP(clk), .CD(n1509), .Q(f42[12]) );
  CFD2QXL \f42_reg[11]  ( .D(s42[11]), .CP(clk), .CD(n1508), .Q(f42[11]) );
  CFD2QXL \f42_reg[10]  ( .D(s42[10]), .CP(clk), .CD(n1491), .Q(f42[10]) );
  CFD2QXL \f42_reg[9]  ( .D(s42[9]), .CP(clk), .CD(n1493), .Q(f42[9]) );
  CFD2QXL \f42_reg[8]  ( .D(s42[8]), .CP(clk), .CD(n1494), .Q(f42[8]) );
  CFD2QXL \f42_reg[7]  ( .D(s42[7]), .CP(clk), .CD(n1496), .Q(f42[7]) );
  CFD2QXL \f42_reg[6]  ( .D(s42[6]), .CP(clk), .CD(n1498), .Q(f42[6]) );
  CFD2QXL \f42_reg[5]  ( .D(s42[5]), .CP(clk), .CD(n1499), .Q(f42[5]) );
  CFD2QXL \f42_reg[4]  ( .D(s42[4]), .CP(clk), .CD(n1501), .Q(f42[4]) );
  CFD2QXL \f42_reg[3]  ( .D(s42[3]), .CP(clk), .CD(n1436), .Q(f42[3]) );
  CFD2QXL \f42_reg[2]  ( .D(s42[2]), .CP(clk), .CD(n1437), .Q(f42[2]) );
  CFD2QXL \f42_reg[1]  ( .D(s42[1]), .CP(clk), .CD(n1439), .Q(f42[1]) );
  CFD2QXL \f52_reg[31]  ( .D(n408), .CP(clk), .CD(n1479), .Q(f52[31]) );
  CFD2QXL \f52_reg[30]  ( .D(n344), .CP(clk), .CD(n1480), .Q(f52[30]) );
  CFD2QXL \f52_reg[29]  ( .D(n410), .CP(clk), .CD(n1482), .Q(f52[29]) );
  CFD2QXL \f52_reg[28]  ( .D(n412), .CP(clk), .CD(n1483), .Q(f52[28]) );
  CFD2QXL \f52_reg[27]  ( .D(n400), .CP(clk), .CD(n1485), .Q(f52[27]) );
  CFD2QXL \f52_reg[26]  ( .D(n402), .CP(clk), .CD(n1487), .Q(f52[26]) );
  CFD2QXL \f52_reg[25]  ( .D(n346), .CP(clk), .CD(n1488), .Q(f52[25]) );
  CFD2QXL \f52_reg[24]  ( .D(n404), .CP(clk), .CD(n1468), .Q(f52[24]) );
  CFD2QXL \f52_reg[23]  ( .D(n406), .CP(clk), .CD(n1469), .Q(f52[23]) );
  CFD2QXL \f52_reg[22]  ( .D(n392), .CP(clk), .CD(n1471), .Q(f52[22]) );
  CFD2QXL \f52_reg[21]  ( .D(n394), .CP(clk), .CD(n1473), .Q(f52[21]) );
  CFD2QXL \f52_reg[20]  ( .D(n348), .CP(clk), .CD(n1474), .Q(f52[20]) );
  CFD2QXL \f52_reg[19]  ( .D(n396), .CP(clk), .CD(n1476), .Q(f52[19]) );
  CFD2QXL \f52_reg[18]  ( .D(n398), .CP(clk), .CD(n1477), .Q(f52[18]) );
  CFD2QXL \f52_reg[17]  ( .D(n384), .CP(clk), .CD(n1501), .Q(f52[17]) );
  CFD2QXL \f52_reg[16]  ( .D(n386), .CP(clk), .CD(n1502), .Q(f52[16]) );
  CFD2QXL \f52_reg[15]  ( .D(n350), .CP(clk), .CD(n1504), .Q(f52[15]) );
  CFD2QXL \f52_reg[14]  ( .D(n388), .CP(clk), .CD(n1505), .Q(f52[14]) );
  CFD2QXL \f52_reg[13]  ( .D(n390), .CP(clk), .CD(n1507), .Q(f52[13]) );
  CFD2QXL \f52_reg[12]  ( .D(n376), .CP(clk), .CD(n1509), .Q(f52[12]) );
  CFD2QXL \f52_reg[11]  ( .D(n378), .CP(clk), .CD(n1510), .Q(f52[11]) );
  CFD2QXL \f52_reg[10]  ( .D(n352), .CP(clk), .CD(n1491), .Q(f52[10]) );
  CFD2QXL \f52_reg[9]  ( .D(n380), .CP(clk), .CD(n1493), .Q(f52[9]) );
  CFD2QXL \f52_reg[8]  ( .D(n382), .CP(clk), .CD(n1494), .Q(f52[8]) );
  CFD2QXL \f52_reg[7]  ( .D(n368), .CP(clk), .CD(n1496), .Q(f52[7]) );
  CFD2QXL \f52_reg[6]  ( .D(n370), .CP(clk), .CD(n1497), .Q(f52[6]) );
  CFD2QXL \f52_reg[5]  ( .D(n354), .CP(clk), .CD(n1499), .Q(f52[5]) );
  CFD2QXL \f52_reg[4]  ( .D(n372), .CP(clk), .CD(n1501), .Q(f52[4]) );
  CFD2QXL \f52_reg[3]  ( .D(n374), .CP(clk), .CD(n1436), .Q(f52[3]) );
  CFD2QXL \f52_reg[2]  ( .D(n364), .CP(clk), .CD(n1437), .Q(f52[2]) );
  CFD2QXL \f52_reg[1]  ( .D(n366), .CP(clk), .CD(n1439), .Q(f52[1]) );
  CFD2QXL \f52_reg[0]  ( .D(n356), .CP(clk), .CD(n1440), .Q(f52[0]) );
  CFD2QXL \f54_reg[29]  ( .D(s54[29]), .CP(clk), .CD(n1483), .Q(f54[29]) );
  CFD2QXL \f54_reg[28]  ( .D(s54[28]), .CP(clk), .CD(n1484), .Q(f54[28]) );
  CFD2QXL \f54_reg[27]  ( .D(s54[27]), .CP(clk), .CD(n1486), .Q(f54[27]) );
  CFD2QXL \f54_reg[26]  ( .D(s54[26]), .CP(clk), .CD(n1488), .Q(f54[26]) );
  CFD2QXL \f54_reg[25]  ( .D(s54[25]), .CP(clk), .CD(n1489), .Q(f54[25]) );
  CFD2QXL \f54_reg[24]  ( .D(s54[24]), .CP(clk), .CD(n1469), .Q(f54[24]) );
  CFD2QXL \f54_reg[23]  ( .D(s54[23]), .CP(clk), .CD(n1470), .Q(f54[23]) );
  CFD2QXL \f54_reg[22]  ( .D(s54[22]), .CP(clk), .CD(n1472), .Q(f54[22]) );
  CFD2QXL \f54_reg[21]  ( .D(s54[21]), .CP(clk), .CD(n1473), .Q(f54[21]) );
  CFD2QXL \f54_reg[20]  ( .D(s54[20]), .CP(clk), .CD(n1475), .Q(f54[20]) );
  CFD2QXL \f54_reg[19]  ( .D(s54[19]), .CP(clk), .CD(n1477), .Q(f54[19]) );
  CFD2QXL \f54_reg[18]  ( .D(s54[18]), .CP(clk), .CD(n1478), .Q(f54[18]) );
  CFD2QXL \f54_reg[17]  ( .D(s54[17]), .CP(clk), .CD(n1502), .Q(f54[17]) );
  CFD2QXL \f54_reg[16]  ( .D(s54[16]), .CP(clk), .CD(n1503), .Q(f54[16]) );
  CFD2QXL \f54_reg[15]  ( .D(s54[15]), .CP(clk), .CD(n1505), .Q(f54[15]) );
  CFD2QXL \f54_reg[14]  ( .D(s54[14]), .CP(clk), .CD(n1507), .Q(f54[14]) );
  CFD2QXL \f54_reg[13]  ( .D(s54[13]), .CP(clk), .CD(n1508), .Q(f54[13]) );
  CFD2QXL \f54_reg[12]  ( .D(s54[12]), .CP(clk), .CD(n1509), .Q(f54[12]) );
  CFD2QXL \f54_reg[11]  ( .D(s54[11]), .CP(clk), .CD(n1490), .Q(f54[11]) );
  CFD2QXL \f54_reg[10]  ( .D(s54[10]), .CP(clk), .CD(n1492), .Q(f54[10]) );
  CFD2QXL \f54_reg[9]  ( .D(s54[9]), .CP(clk), .CD(n1494), .Q(f54[9]) );
  CFD2QXL \f54_reg[8]  ( .D(s54[8]), .CP(clk), .CD(n1495), .Q(f54[8]) );
  CFD2QXL \f54_reg[7]  ( .D(s54[7]), .CP(clk), .CD(n1497), .Q(f54[7]) );
  CFD2QXL \f54_reg[6]  ( .D(s54[6]), .CP(clk), .CD(n1498), .Q(f54[6]) );
  CFD2QXL \f54_reg[5]  ( .D(s54[5]), .CP(clk), .CD(n1500), .Q(f54[5]) );
  CFD2QXL \f54_reg[4]  ( .D(s54[4]), .CP(clk), .CD(n1435), .Q(f54[4]) );
  CFD2QXL \f54_reg[3]  ( .D(s54[3]), .CP(clk), .CD(n1437), .Q(f54[3]) );
  CFD2QXL \f54_reg[2]  ( .D(s54[2]), .CP(clk), .CD(n1438), .Q(f54[2]) );
  CFD2QXL \f61_reg[29]  ( .D(s61[29]), .CP(clk), .CD(n1482), .Q(f61[29]) );
  CFD2QXL \f61_reg[28]  ( .D(s61[28]), .CP(clk), .CD(n1484), .Q(f61[28]) );
  CFD2QXL \f61_reg[27]  ( .D(s61[27]), .CP(clk), .CD(n1486), .Q(f61[27]) );
  CFD2QXL \f61_reg[26]  ( .D(s61[26]), .CP(clk), .CD(n1487), .Q(f61[26]) );
  CFD2QXL \f61_reg[25]  ( .D(s61[25]), .CP(clk), .CD(n1489), .Q(f61[25]) );
  CFD2QXL \f61_reg[24]  ( .D(s61[24]), .CP(clk), .CD(n1468), .Q(f61[24]) );
  CFD2QXL \f61_reg[23]  ( .D(s61[23]), .CP(clk), .CD(n1470), .Q(f61[23]) );
  CFD2QXL \f61_reg[22]  ( .D(s61[22]), .CP(clk), .CD(n1471), .Q(f61[22]) );
  CFD2QXL \f61_reg[21]  ( .D(s61[21]), .CP(clk), .CD(n1473), .Q(f61[21]) );
  CFD2QXL \f61_reg[20]  ( .D(s61[20]), .CP(clk), .CD(n1475), .Q(f61[20]) );
  CFD2QXL \f61_reg[19]  ( .D(s61[19]), .CP(clk), .CD(n1476), .Q(f61[19]) );
  CFD2QXL \f61_reg[18]  ( .D(s61[18]), .CP(clk), .CD(n1478), .Q(f61[18]) );
  CFD2QXL \f61_reg[17]  ( .D(s61[17]), .CP(clk), .CD(n1501), .Q(f61[17]) );
  CFD2QXL \f61_reg[16]  ( .D(s61[16]), .CP(clk), .CD(n1503), .Q(f61[16]) );
  CFD2QXL \f61_reg[15]  ( .D(s61[15]), .CP(clk), .CD(n1504), .Q(f61[15]) );
  CFD2QXL \f61_reg[14]  ( .D(s61[14]), .CP(clk), .CD(n1506), .Q(f61[14]) );
  CFD2QXL \f61_reg[13]  ( .D(s61[13]), .CP(clk), .CD(n1507), .Q(f61[13]) );
  CFD2QXL \f61_reg[12]  ( .D(s61[12]), .CP(clk), .CD(n1508), .Q(f61[12]) );
  CFD2QXL \f61_reg[11]  ( .D(s61[11]), .CP(clk), .CD(n1490), .Q(f61[11]) );
  CFD2QXL \f61_reg[10]  ( .D(s61[10]), .CP(clk), .CD(n1492), .Q(f61[10]) );
  CFD2QXL \f61_reg[9]  ( .D(s61[9]), .CP(clk), .CD(n1493), .Q(f61[9]) );
  CFD2QXL \f61_reg[8]  ( .D(s61[8]), .CP(clk), .CD(n1495), .Q(f61[8]) );
  CFD2QXL \f61_reg[7]  ( .D(s61[7]), .CP(clk), .CD(n1496), .Q(f61[7]) );
  CFD2QXL \f61_reg[6]  ( .D(s61[6]), .CP(clk), .CD(n1498), .Q(f61[6]) );
  CFD2QXL \f61_reg[5]  ( .D(s61[5]), .CP(clk), .CD(n1500), .Q(f61[5]) );
  CFD2QXL \f61_reg[4]  ( .D(s61[4]), .CP(clk), .CD(n1435), .Q(f61[4]) );
  CFD2QXL \f61_reg[3]  ( .D(s61[3]), .CP(clk), .CD(n1436), .Q(f61[3]) );
  CFD2QXL \f61_reg[2]  ( .D(s61[2]), .CP(clk), .CD(n1438), .Q(f61[2]) );
  CFD2QXL \f61_reg[1]  ( .D(s61[1]), .CP(clk), .CD(n1439), .Q(f61[1]) );
  CFD2QXL pushOut_reg ( .D(n561), .CP(clk), .CD(n1463), .Q(pushZ) );
  CFD2QXL \res_reg[0]  ( .D(n563), .CP(clk), .CD(n1440), .Q(Z[0]) );
  CFD2QXL \res_reg[1]  ( .D(n564), .CP(clk), .CD(n1439), .Q(Z[1]) );
  CFD2QXL \res_reg[2]  ( .D(n307), .CP(clk), .CD(n1437), .Q(Z[2]) );
  CFD2QXL \res_reg[3]  ( .D(n565), .CP(clk), .CD(n1436), .Q(Z[3]) );
  CFD2QXL \res_reg[4]  ( .D(n557), .CP(clk), .CD(n1500), .Q(Z[4]) );
  CFD2QXL \res_reg[5]  ( .D(n558), .CP(clk), .CD(n1499), .Q(Z[5]) );
  CFD2QXL \res_reg[6]  ( .D(n559), .CP(clk), .CD(n1497), .Q(Z[6]) );
  CFD2QXL \res_reg[7]  ( .D(n308), .CP(clk), .CD(n1496), .Q(Z[7]) );
  CFD2QXL \res_reg[8]  ( .D(n560), .CP(clk), .CD(n1494), .Q(Z[8]) );
  CFD2QXL \res_reg[9]  ( .D(n553), .CP(clk), .CD(n1492), .Q(Z[9]) );
  CFD2QXL \res_reg[10]  ( .D(n554), .CP(clk), .CD(n1491), .Q(Z[10]) );
  CFD2QXL \res_reg[11]  ( .D(n555), .CP(clk), .CD(n1509), .Q(Z[11]) );
  CFD2QXL \res_reg[12]  ( .D(n309), .CP(clk), .CD(n1509), .Q(Z[12]) );
  CFD2QXL \res_reg[13]  ( .D(n556), .CP(clk), .CD(n1507), .Q(Z[13]) );
  CFD2QXL \res_reg[14]  ( .D(n549), .CP(clk), .CD(n1505), .Q(Z[14]) );
  CFD2QXL \res_reg[15]  ( .D(n550), .CP(clk), .CD(n1504), .Q(Z[15]) );
  CFD2QXL \res_reg[16]  ( .D(n551), .CP(clk), .CD(n1502), .Q(Z[16]) );
  CFD2QXL \res_reg[17]  ( .D(n310), .CP(clk), .CD(n1479), .Q(Z[17]) );
  CFD2QXL \res_reg[18]  ( .D(n552), .CP(clk), .CD(n1477), .Q(Z[18]) );
  CFD2QXL \res_reg[19]  ( .D(n545), .CP(clk), .CD(n1476), .Q(Z[19]) );
  CFD2QXL \res_reg[20]  ( .D(n546), .CP(clk), .CD(n1474), .Q(Z[20]) );
  CFD2QXL \res_reg[21]  ( .D(n547), .CP(clk), .CD(n1472), .Q(Z[21]) );
  CFD2QXL \res_reg[22]  ( .D(n311), .CP(clk), .CD(n1471), .Q(Z[22]) );
  CFD2QXL \res_reg[23]  ( .D(n548), .CP(clk), .CD(n1469), .Q(Z[23]) );
  CFD2QXL \res_reg[24]  ( .D(n541), .CP(clk), .CD(n1473), .Q(Z[24]) );
  CFD2QXL \res_reg[25]  ( .D(n542), .CP(clk), .CD(n1488), .Q(Z[25]) );
  CFD2QXL \res_reg[26]  ( .D(n543), .CP(clk), .CD(n1487), .Q(Z[26]) );
  CFD2QXL \res_reg[27]  ( .D(n312), .CP(clk), .CD(n1485), .Q(Z[27]) );
  CFD2QXL \res_reg[28]  ( .D(n544), .CP(clk), .CD(n1483), .Q(Z[28]) );
  CFD2QXL \res_reg[29]  ( .D(n538), .CP(clk), .CD(n1482), .Q(Z[29]) );
  CFD2QXL \res_reg[30]  ( .D(n539), .CP(clk), .CD(n1480), .Q(Z[30]) );
  CFD2QXL \res_reg[31]  ( .D(n540), .CP(clk), .CD(n1424), .Q(Z[31]) );
  CFD2QXL \f21_reg[10]  ( .D(n189), .CP(clk), .CD(n1434), .Q(f21[10]) );
  CFD2QXL \f21_reg[9]  ( .D(n190), .CP(clk), .CD(n1457), .Q(f21[9]) );
  CFD2QXL \f01_reg[16]  ( .D(n528), .CP(clk), .CD(n1431), .Q(f01[16]) );
  CFD2QXL \f01_reg[4]  ( .D(n522), .CP(clk), .CD(n1460), .Q(f01[4]) );
  CFD2QX1 \f14_reg[21]  ( .D(w2[21]), .CP(clk), .CD(n1475), .Q(f14[21]) );
  CFD2QX1 \f36_reg[7]  ( .D(n265), .CP(clk), .CD(n1458), .Q(f36[7]) );
  CFD2QX1 \f14_reg[17]  ( .D(w2[17]), .CP(clk), .CD(n1504), .Q(f14[17]) );
  CFD2QX1 \f21_reg[4]  ( .D(n183), .CP(clk), .CD(n1460), .Q(f21[4]) );
  CFD2QX1 \f21_reg[3]  ( .D(n262), .CP(clk), .CD(n1461), .Q(f21[3]) );
  CFD2QX1 \f21_reg[5]  ( .D(n185), .CP(clk), .CD(n1459), .Q(f21[5]) );
  CFD2QX1 \f14_reg[13]  ( .D(w2[13]), .CP(clk), .CD(n1510), .Q(f14[13]) );
  CFD2QX1 \f14_reg[11]  ( .D(w2[11]), .CP(clk), .CD(n1492), .Q(f14[11]) );
  CFD2QX1 \f14_reg[19]  ( .D(w2[19]), .CP(clk), .CD(n1478), .Q(f14[19]) );
  CFD2QX1 \f14_reg[15]  ( .D(w2[15]), .CP(clk), .CD(n1507), .Q(f14[15]) );
  CFD2QX1 \f01_reg[11]  ( .D(n250), .CP(clk), .CD(n1434), .Q(f01[11]) );
  CFD2QX1 \captA_reg[20]  ( .D(n170), .CP(clk), .CD(n1428), .Q(captA[20]) );
  CFD2QX1 \captA_reg[19]  ( .D(n169), .CP(clk), .CD(n1429), .Q(captA[19]) );
  CFD2QX1 \captA_reg[18]  ( .D(n168), .CP(clk), .CD(n1429), .Q(captA[18]) );
  CFD2QX1 \captA_reg[16]  ( .D(n166), .CP(clk), .CD(n1431), .Q(captA[16]) );
  CFD2QX1 \f03_reg[1]  ( .D(n249), .CP(clk), .CD(n1456), .Q(f03[1]) );
  CFD2QX1 \captC_reg[20]  ( .D(n106), .CP(clk), .CD(n1447), .Q(captC[20]) );
  CFD2QX1 \captB_reg[20]  ( .D(n138), .CP(clk), .CD(n1475), .Q(captB[20]) );
  CFD2QX1 \captB_reg[19]  ( .D(n137), .CP(clk), .CD(n1477), .Q(captB[19]) );
  CFD2QX1 \captC_reg[19]  ( .D(n105), .CP(clk), .CD(n1448), .Q(captC[19]) );
  CFD2QX1 \captB_reg[18]  ( .D(n136), .CP(clk), .CD(n1479), .Q(captB[18]) );
  CFD2QX1 \captC_reg[18]  ( .D(n104), .CP(clk), .CD(n1448), .Q(captC[18]) );
  CFD2QX1 \captB_reg[16]  ( .D(n134), .CP(clk), .CD(n1504), .Q(captB[16]) );
  CFD2QX1 \captC_reg[16]  ( .D(n102), .CP(clk), .CD(n1449), .Q(captC[16]) );
  CFD2QX1 \captA_reg[15]  ( .D(n165), .CP(clk), .CD(n1431), .Q(captA[15]) );
  CFD2QX1 \captA_reg[14]  ( .D(n164), .CP(clk), .CD(n1432), .Q(captA[14]) );
  CFD2QX1 \captA_reg[13]  ( .D(n163), .CP(clk), .CD(n1433), .Q(captA[13]) );
  CFD2QX1 \captB_reg[13]  ( .D(n131), .CP(clk), .CD(n1508), .Q(captB[13]) );
  CFD2QX1 \captA_reg[12]  ( .D(n162), .CP(clk), .CD(n1433), .Q(captA[12]) );
  CFD2QX1 \captA_reg[11]  ( .D(n161), .CP(clk), .CD(n1434), .Q(captA[11]) );
  CFD2QX1 \captC_reg[11]  ( .D(n97), .CP(clk), .CD(n1451), .Q(captC[11]) );
  CFD2QX2 \captB_reg[3]  ( .D(n121), .CP(clk), .CD(n1437), .Q(captB[3]) );
  CFD2QX1 \captB_reg[11]  ( .D(n129), .CP(clk), .CD(n1491), .Q(captB[11]) );
  CFD2QX1 \captB_reg[14]  ( .D(n132), .CP(clk), .CD(n1507), .Q(captB[14]) );
  CFD2QX1 \captB_reg[15]  ( .D(n133), .CP(clk), .CD(n1505), .Q(captB[15]) );
  CFD2QX1 \captC_reg[15]  ( .D(n101), .CP(clk), .CD(n1450), .Q(captC[15]) );
  CFD2QX1 \captC_reg[13]  ( .D(n99), .CP(clk), .CD(n1450), .Q(captC[13]) );
  CFD2QX1 \captC_reg[12]  ( .D(n98), .CP(clk), .CD(n1451), .Q(captC[12]) );
  CFD2QX1 \captB_reg[12]  ( .D(n130), .CP(clk), .CD(n1510), .Q(captB[12]) );
  CFD2QX2 \captC_reg[4]  ( .D(n90), .CP(clk), .CD(n1455), .Q(captC[4]) );
  CFD2QX2 \captA_reg[3]  ( .D(n153), .CP(clk), .CD(n1461), .Q(captA[3]) );
  CFD2QX2 \captC_reg[3]  ( .D(n89), .CP(clk), .CD(n1455), .Q(captC[3]) );
  CFD2QX2 \captB_reg[0]  ( .D(n118), .CP(clk), .CD(n1442), .Q(captB[0]) );
  CFD2QX1 \f12_reg[26]  ( .D(w1[26]), .CP(clk), .CD(n1424), .Q(f12[26]) );
  CFD2QX1 \f02_reg[26]  ( .D(n313), .CP(clk), .CD(n1488), .Q(f02[26]) );
  CFD2QX2 \f02_reg[24]  ( .D(n513), .CP(clk), .CD(n1469), .Q(f02[24]) );
  CFD2QX1 \f11_reg[18]  ( .D(f01[18]), .CP(clk), .CD(n1429), .Q(f11[18]) );
  CFD2QX1 \f11_reg[16]  ( .D(f01[16]), .CP(clk), .CD(n1430), .Q(f11[16]) );
  CFD2QX1 \f03_reg[23]  ( .D(n512), .CP(clk), .CD(n1451), .Q(f03[23]) );
  CFD2QX2 \f02_reg[23]  ( .D(n273), .CP(clk), .CD(n1470), .Q(f02[23]) );
  CFD2QXL \f21_reg[6]  ( .D(n274), .CP(clk), .CD(n1459), .Q(f21[6]) );
  CFD2QXL \f01_reg[17]  ( .D(n279), .CP(clk), .CD(n1430), .Q(f01[17]) );
  CFD2QXL \f14_reg[25]  ( .D(w2[25]), .CP(clk), .CD(n1469), .Q(f14[25]) );
  CFD2QXL \f14_reg[23]  ( .D(w2[23]), .CP(clk), .CD(n1472), .Q(f14[23]) );
  CFD2QXL \f36_reg[12]  ( .D(n282), .CP(clk), .CD(n1433), .Q(f36[12]) );
  CFD2QXL \f36_reg[13]  ( .D(n280), .CP(clk), .CD(n1432), .Q(f36[13]) );
  CFD2QXL \f14_reg[14]  ( .D(w2[14]), .CP(clk), .CD(n1508), .Q(f14[14]) );
  CFD2QXL \f14_reg[0]  ( .D(w2[0]), .CP(clk), .CD(n1442), .Q(f14[0]) );
  CFD2QX2 \captC_reg[0]  ( .D(n86), .CP(clk), .CD(n1457), .Q(captC[0]) );
  CFD2QX2 \captA_reg[0]  ( .D(n150), .CP(clk), .CD(n1463), .Q(captA[0]) );
  CFD2QX2 \captA_reg[8]  ( .D(n158), .CP(clk), .CD(n1458), .Q(captA[8]) );
  CFD2QX2 \captB_reg[8]  ( .D(n126), .CP(clk), .CD(n1496), .Q(captB[8]) );
  CFD2QX2 \captA_reg[7]  ( .D(n157), .CP(clk), .CD(n1458), .Q(captA[7]) );
  CFD2QX2 \captB_reg[7]  ( .D(n125), .CP(clk), .CD(n1497), .Q(captB[7]) );
  CFD2QX2 \captA_reg[5]  ( .D(n155), .CP(clk), .CD(n1460), .Q(captA[5]) );
  CFD2QX2 \captB_reg[4]  ( .D(n122), .CP(clk), .CD(n1435), .Q(captB[4]) );
  CFD2QX2 \captA_reg[4]  ( .D(n154), .CP(clk), .CD(n1460), .Q(captA[4]) );
  CFD2QX2 \captC_reg[8]  ( .D(n94), .CP(clk), .CD(n1453), .Q(captC[8]) );
  CFD2QX2 \captC_reg[6]  ( .D(n92), .CP(clk), .CD(n1454), .Q(captC[6]) );
  CFD2QX2 \captC_reg[7]  ( .D(n93), .CP(clk), .CD(n1453), .Q(captC[7]) );
  CFD2QX2 \captC_reg[5]  ( .D(n91), .CP(clk), .CD(n1454), .Q(captC[5]) );
  CFD2QX2 \captB_reg[5]  ( .D(n123), .CP(clk), .CD(n1500), .Q(captB[5]) );
  CFD2QXL \f14_reg[12]  ( .D(w2[12]), .CP(clk), .CD(n1491), .Q(f14[12]) );
  CFD2QXL \f03_reg[25]  ( .D(n220), .CP(clk), .CD(n1467), .Q(f03[25]) );
  CFD2QXL \f03_reg[24]  ( .D(n222), .CP(clk), .CD(n1467), .Q(f03[24]) );
  CFD2QX4 \f03_reg[9]  ( .D(n224), .CP(clk), .CD(n1452), .Q(f03[9]) );
  CFD2QX1 \captA_reg[10]  ( .D(n160), .CP(clk), .CD(n1435), .Q(captA[10]) );
  CFD2QX1 \captA_reg[9]  ( .D(n159), .CP(clk), .CD(n1457), .Q(captA[9]) );
  CFD2QX1 \captB_reg[9]  ( .D(n127), .CP(clk), .CD(n1494), .Q(captB[9]) );
  CFD2QX1 \captC_reg[9]  ( .D(n95), .CP(clk), .CD(n1452), .Q(captC[9]) );
  CFD2QX1 \f36_reg[5]  ( .D(n358), .CP(clk), .CD(n1459), .Q(f36[5]) );
  CFD2QX2 \f03_reg[11]  ( .D(n509), .CP(clk), .CD(n1451), .Q(f03[11]) );
  CFD2QX1 \f01_reg[23]  ( .D(n361), .CP(clk), .CD(n1426), .Q(f01[23]) );
  CFD2QX4 \f02_reg[21]  ( .D(n459), .CP(clk), .CD(n1474), .Q(f02[21]) );
  CFD2QX1 \captC_reg[10]  ( .D(n96), .CP(clk), .CD(n1452), .Q(captC[10]) );
  CFD2QX1 \captB_reg[10]  ( .D(n128), .CP(clk), .CD(n1492), .Q(captB[10]) );
  CFD2QXL \f14_reg[9]  ( .D(w2[9]), .CP(clk), .CD(n1496), .Q(f14[9]) );
  CFD2QXL \f14_reg[5]  ( .D(w2[5]), .CP(clk), .CD(n1435), .Q(f14[5]) );
  CFD2QXL \f14_reg[3]  ( .D(w2[3]), .CP(clk), .CD(n1438), .Q(f14[3]) );
  CFD2QXL \f01_reg[15]  ( .D(n505), .CP(clk), .CD(n1431), .Q(f01[15]) );
  CFD2QXL \f01_reg[13]  ( .D(n507), .CP(clk), .CD(n1432), .Q(f01[13]) );
  CFD2QX1 \f02_reg[3]  ( .D(n203), .CP(clk), .CD(n1437), .Q(f02[3]) );
  CFD2QX1 \f12_reg[24]  ( .D(w1[24]), .CP(clk), .CD(n1426), .Q(f12[24]) );
  CFD2QX2 \f12_reg[22]  ( .D(w1[22]), .CP(clk), .CD(n1428), .Q(f12[22]) );
  CFD2QX4 \f03_reg[7]  ( .D(n204), .CP(clk), .CD(n1453), .Q(f03[7]) );
  CFD2QX1 \f01_reg[29]  ( .D(n205), .CP(clk), .CD(n1444), .Q(f01[29]) );
  CFD2QX1 \f03_reg[22]  ( .D(n206), .CP(clk), .CD(n1446), .Q(f03[22]) );
  CFD2QX4 \f03_reg[6]  ( .D(n208), .CP(clk), .CD(n1453), .Q(f03[6]) );
  CFD2QX4 \f03_reg[8]  ( .D(n207), .CP(clk), .CD(n1452), .Q(f03[8]) );
  CFD2QX1 \f02_reg[4]  ( .D(n209), .CP(clk), .CD(n1435), .Q(f02[4]) );
  CFD2XL \f53_reg[31]  ( .D(w11[31]), .CP(clk), .CD(n1442), .Q(n1420) );
  CFD2QX1 \f02_reg[13]  ( .D(n501), .CP(clk), .CD(n1509), .Q(f02[13]) );
  CFD2QX1 \f01_reg[5]  ( .D(n499), .CP(clk), .CD(n1460), .Q(f01[5]) );
  CFD2QX1 \f02_reg[1]  ( .D(n314), .CP(clk), .CD(n1440), .Q(f02[1]) );
  CFD2QX1 \f11_reg[3]  ( .D(n315), .CP(clk), .CD(n1461), .Q(f11[3]) );
  CFD2QX1 \f12_reg[28]  ( .D(w1[28]), .CP(clk), .CD(n1445), .Q(f12[28]) );
  CFD2QX1 \f11_reg[19]  ( .D(n493), .CP(clk), .CD(n1428), .Q(f11[19]) );
  CFD2QX1 \f01_reg[19]  ( .D(n496), .CP(clk), .CD(n1428), .Q(f01[19]) );
  CFD2QX1 \f02_reg[9]  ( .D(n318), .CP(clk), .CD(n1494), .Q(f02[9]) );
  CFD2QX1 \f02_reg[8]  ( .D(n491), .CP(clk), .CD(n1495), .Q(f02[8]) );
  CFD2QX1 \f01_reg[7]  ( .D(n485), .CP(clk), .CD(n1458), .Q(f01[7]) );
  CFD2QX1 \f01_reg[0]  ( .D(n484), .CP(clk), .CD(n1463), .Q(f01[0]) );
  CFD2QX1 \f01_reg[1]  ( .D(n482), .CP(clk), .CD(n1462), .Q(f01[1]) );
  CFD2QX1 \f14_reg[7]  ( .D(w2[7]), .CP(clk), .CD(n1499), .Q(f14[7]) );
  CFD2QX1 \f11_reg[21]  ( .D(n438), .CP(clk), .CD(n1427), .Q(f11[21]) );
  CFD2QX1 \f01_reg[21]  ( .D(n441), .CP(clk), .CD(n1427), .Q(f01[21]) );
  CFD2QX2 \captC_reg[2]  ( .D(n88), .CP(clk), .CD(n1456), .Q(captC[2]) );
  CFD2QX1 \f03_reg[2]  ( .D(n480), .CP(clk), .CD(n1455), .Q(f03[2]) );
  CFD2QX2 \f01_reg[2]  ( .D(n442), .CP(clk), .CD(n1462), .Q(f01[2]) );
  CFD2QX1 \f01_reg[12]  ( .D(n335), .CP(clk), .CD(n1433), .Q(f01[12]) );
  CFD2QX1 \f11_reg[12]  ( .D(n444), .CP(clk), .CD(n1433), .Q(f11[12]) );
  CFD2QX1 \f12_reg[25]  ( .D(w1[25]), .CP(clk), .CD(n1425), .Q(f12[25]) );
  CFD2QX2 \captB_reg[2]  ( .D(n120), .CP(clk), .CD(n1439), .Q(captB[2]) );
  CFD2QX4 \f02_reg[2]  ( .D(n271), .CP(clk), .CD(n1438), .Q(f02[2]) );
  CFD2QX1 \f11_reg[1]  ( .D(n210), .CP(clk), .CD(n1462), .Q(f11[1]) );
  CFD2QX1 \f36_reg[0]  ( .D(n215), .CP(clk), .CD(n1463), .Q(f36[0]) );
  CFD2QX2 \f11_reg[20]  ( .D(n218), .CP(clk), .CD(n1428), .Q(f11[20]) );
  CFD2QX1 \f01_reg[20]  ( .D(n213), .CP(clk), .CD(n1428), .Q(f01[20]) );
  CFD2XL \f32_reg[31]  ( .D(w8[31]), .CP(clk), .CD(n1479), .Q(n1419) );
  CFD2XL \f31_reg[30]  ( .D(w7[30]), .CP(clk), .CD(n1481), .Q(n1418) );
  CFD2QX1 \f11_reg[2]  ( .D(n479), .CP(clk), .CD(n1461), .Q(f11[2]) );
  CFD2QX1 \f36_reg[2]  ( .D(n257), .CP(clk), .CD(n1461), .Q(f36[2]) );
  CFD2QX1 \f21_reg[2]  ( .D(n254), .CP(clk), .CD(n1461), .Q(f21[2]) );
  CFD2QX1 \f11_reg[22]  ( .D(f01[22]), .CP(clk), .CD(n1427), .Q(f11[22]) );
  CFD2X1 \f36_reg[1]  ( .D(n473), .CP(clk), .CD(n1462), .Q(f36[1]) );
  CFD2QX1 \f21_reg[1]  ( .D(n251), .CP(clk), .CD(n1462), .Q(f21[1]) );
  CFD2QX2 \f11_reg[0]  ( .D(n471), .CP(clk), .CD(n1463), .Q(f11[0]) );
  CFD2QX1 \f21_reg[0]  ( .D(n468), .CP(clk), .CD(n1463), .Q(f21[0]) );
  CFD2QXL \f32_reg[30]  ( .D(w8[30]), .CP(clk), .CD(n1480), .Q(f32[30]) );
  CFD2QX1 \f01_reg[6]  ( .D(n457), .CP(clk), .CD(n1459), .Q(f01[6]) );
  CFD2QX1 \f11_reg[6]  ( .D(n456), .CP(clk), .CD(n1459), .Q(f11[6]) );
  CFD2QX1 \f36_reg[4]  ( .D(n449), .CP(clk), .CD(n1460), .Q(f36[4]) );
  CFD2QX2 \f01_reg[8]  ( .D(n454), .CP(clk), .CD(n1458), .Q(f01[8]) );
  CFD2QX1 \f01_reg[9]  ( .D(n452), .CP(clk), .CD(n1457), .Q(f01[9]) );
  CFD2QX1 \f02_reg[6]  ( .D(n447), .CP(clk), .CD(n1499), .Q(f02[6]) );
  CFD2QX1 \f13_reg[6]  ( .D(n445), .CP(clk), .CD(n1498), .Q(f13[6]) );
  CFD2QX4 \f03_reg[17]  ( .D(n330), .CP(clk), .CD(n1448), .Q(f03[17]) );
  CFD2QX2 \f11_reg[17]  ( .D(n333), .CP(clk), .CD(n1430), .Q(f11[17]) );
  CFD2QX1 \f36_reg[3]  ( .D(n327), .CP(clk), .CD(n1461), .Q(f36[3]) );
  CFD2QX1 \f11_reg[7]  ( .D(n321), .CP(clk), .CD(n1458), .Q(f11[7]) );
  CFD2QX1 \f01_reg[14]  ( .D(n324), .CP(clk), .CD(n1432), .Q(f01[14]) );
  CFD2QX1 \f11_reg[14]  ( .D(n184), .CP(clk), .CD(n1432), .Q(f11[14]) );
  CFD2QX2 \captC_reg[14]  ( .D(n100), .CP(clk), .CD(n1513), .Q(captC[14]) );
  CFD2QX1 \f11_reg[25]  ( .D(n769), .CP(clk), .CD(n1424), .Q(f11[25]) );
  CFD2QX2 \f11_reg[8]  ( .D(n808), .CP(clk), .CD(n1457), .Q(f11[8]) );
  CFD2QX1 \f11_reg[9]  ( .D(n816), .CP(clk), .CD(n1457), .Q(f11[9]) );
  CFD2QX1 \f11_reg[5]  ( .D(n803), .CP(clk), .CD(n1459), .Q(f11[5]) );
  CFD2QX2 \f36_reg[9]  ( .D(n949), .CP(clk), .CD(n1457), .Q(f36[9]) );
  CFD2QX1 \f03_reg[0]  ( .D(n524), .CP(clk), .CD(n1456), .Q(f03[0]) );
  CFD2QX1 \f11_reg[15]  ( .D(n806), .CP(clk), .CD(n1431), .Q(f11[15]) );
  CFD2QX2 \f02_reg[17]  ( .D(n201), .CP(clk), .CD(n1502), .Q(f02[17]) );
  CFD2QX1 \captB_reg[17]  ( .D(n135), .CP(clk), .CD(n1502), .Q(captB[17]) );
  CFD2QX1 \f11_reg[10]  ( .D(n200), .CP(clk), .CD(n1434), .Q(f11[10]) );
  CFD2QX1 \f01_reg[10]  ( .D(n531), .CP(clk), .CD(n1434), .Q(f01[10]) );
  CFD2QX1 \f11_reg[4]  ( .D(n284), .CP(clk), .CD(n1460), .Q(f11[4]) );
  CFD2QX1 \f02_reg[28]  ( .D(n736), .CP(clk), .CD(n1485), .Q(f02[28]) );
  CFD2QX1 \f02_reg[7]  ( .D(n487), .CP(clk), .CD(n1497), .Q(f02[7]) );
  CFD2QX1 \f02_reg[0]  ( .D(n678), .CP(clk), .CD(n1441), .Q(f02[0]) );
  CFD2QX1 \f02_reg[5]  ( .D(n682), .CP(clk), .CD(n1500), .Q(f02[5]) );
  CFD2QX1 \f03_reg[5]  ( .D(n655), .CP(clk), .CD(n1454), .Q(f03[5]) );
  CFD2QX1 \f03_reg[4]  ( .D(n653), .CP(clk), .CD(n1454), .Q(f03[4]) );
  CFD2QX1 \f03_reg[3]  ( .D(n651), .CP(clk), .CD(n1455), .Q(f03[3]) );
  CFD2QX1 \f12_reg[18]  ( .D(w1[18]), .CP(clk), .CD(n1430), .Q(f12[18]) );
  CFD2QX1 \captA_reg[6]  ( .D(n156), .CP(clk), .CD(n1459), .Q(captA[6]) );
  CFD2QX1 \captB_reg[6]  ( .D(n124), .CP(clk), .CD(n1499), .Q(captB[6]) );
  CFD2QXL \f13_reg[8]  ( .D(n489), .CP(clk), .CD(n1494), .Q(f13[8]) );
  CFD2QX1 \captA_reg[2]  ( .D(n152), .CP(clk), .CD(n1462), .Q(captA[2]) );
  CFD2QX1 \captC_reg[17]  ( .D(n103), .CP(clk), .CD(n1449), .Q(captC[17]) );
  CFD2QX2 \f12_reg[5]  ( .D(w1[5]), .CP(clk), .CD(n1511), .Q(f12[5]) );
  CFD2QX1 \f36_reg[8]  ( .D(n947), .CP(clk), .CD(n1457), .Q(f36[8]) );
  CFD2QX4 \f12_reg[2]  ( .D(w1[2]), .CP(clk), .CD(n1462), .Q(f12[2]) );
  CFD2QX1 \f11_reg[13]  ( .D(n810), .CP(clk), .CD(n1432), .Q(f11[13]) );
  CFD2QX2 \f12_reg[23]  ( .D(w1[23]), .CP(clk), .CD(n1511), .Q(f12[23]) );
  CFD2QX1 \f11_reg[24]  ( .D(n773), .CP(clk), .CD(n1425), .Q(f11[24]) );
  CFD2QX1 \f14_reg[2]  ( .D(w2[2]), .CP(clk), .CD(n1440), .Q(f14[2]) );
  CFD2QX4 \f02_reg[12]  ( .D(n686), .CP(clk), .CD(n1510), .Q(f02[12]) );
  CFD2QX2 \captA_reg[17]  ( .D(n167), .CP(clk), .CD(n1430), .Q(captA[17]) );
  CFD2QX4 \f12_reg[10]  ( .D(w1[10]), .CP(clk), .CD(n1457), .Q(f12[10]) );
  CFD2QX1 \captC_reg[22]  ( .D(n108), .CP(clk), .CD(n1446), .Q(captC[22]) );
  CIVX4 U183 ( .A(n187), .Z(n188) );
  CNIVX1 U184 ( .A(n260), .Z(n183) );
  CNIVX1 U185 ( .A(f01[14]), .Z(n184) );
  CNIVX1 U186 ( .A(n466), .Z(n185) );
  CNIVX1 U187 ( .A(f02[21]), .Z(n186) );
  CIVX2 U188 ( .A(n526), .Z(n187) );
  CNIVX1 U189 ( .A(n534), .Z(n189) );
  CNIVX1 U190 ( .A(n536), .Z(n190) );
  CNIVX1 U191 ( .A(n703), .Z(n191) );
  CNIVX1 U192 ( .A(n193), .Z(n192) );
  CNIVX1 U193 ( .A(n194), .Z(n193) );
  CNIVX1 U194 ( .A(f11[25]), .Z(n194) );
  CNIVX1 U195 ( .A(f11[23]), .Z(n195) );
  CNIVX1 U196 ( .A(f11[24]), .Z(n196) );
  CNIVX1 U197 ( .A(n776), .Z(n197) );
  CNIVXL U198 ( .A(f02[28]), .Z(n782) );
  CNIVX1 U199 ( .A(n782), .Z(n198) );
  CNIVX1 U200 ( .A(n819), .Z(n199) );
  CNIVX1 U201 ( .A(f01[10]), .Z(n200) );
  CNIVX1 U202 ( .A(n326), .Z(n201) );
  CNIVX1 U203 ( .A(captB[17]), .Z(n202) );
  CIVX1 U204 ( .A(n1514), .Z(n1515) );
  CIVX4 U205 ( .A(n1422), .Z(n1423) );
  CIVX2 U206 ( .A(w5[22]), .Z(n1422) );
  CNIVX4 U207 ( .A(n526), .Z(n527) );
  CIVX4 U208 ( .A(n502), .Z(n503) );
  CNIVX1 U209 ( .A(n515), .Z(n203) );
  CNIVX1 U210 ( .A(n227), .Z(n204) );
  CNIVX1 U211 ( .A(captA[29]), .Z(n205) );
  CNIVX1 U212 ( .A(captC[22]), .Z(n206) );
  CNIVX1 U213 ( .A(n225), .Z(n207) );
  CNIVX1 U214 ( .A(n226), .Z(n208) );
  CNIVX1 U215 ( .A(n228), .Z(n209) );
  CNIVX1 U216 ( .A(n211), .Z(n210) );
  CNIVX1 U217 ( .A(n212), .Z(n211) );
  CNIVX1 U218 ( .A(f01[1]), .Z(n212) );
  CNIVX1 U219 ( .A(n214), .Z(n213) );
  CNIVX1 U220 ( .A(n248), .Z(n214) );
  CNIVX1 U221 ( .A(n216), .Z(n215) );
  CNIVX1 U222 ( .A(n217), .Z(n216) );
  CNIVX1 U223 ( .A(f21[0]), .Z(n217) );
  CNIVX1 U224 ( .A(n219), .Z(n218) );
  CNIVX1 U225 ( .A(f01[20]), .Z(n219) );
  CNIVX1 U226 ( .A(n221), .Z(n220) );
  CNIVX1 U227 ( .A(captC[25]), .Z(n221) );
  CNIVX1 U228 ( .A(n223), .Z(n222) );
  CNIVX1 U229 ( .A(captC[24]), .Z(n223) );
  CNIVX1 U230 ( .A(n362), .Z(n224) );
  CNIVX1 U231 ( .A(captC[8]), .Z(n225) );
  CNIVX1 U232 ( .A(captC[6]), .Z(n226) );
  CNIVX1 U233 ( .A(captC[7]), .Z(n227) );
  CNIVX1 U234 ( .A(captB[4]), .Z(n228) );
  CNIVX1 U235 ( .A(f02[12]), .Z(n229) );
  CNIVX1 U236 ( .A(n231), .Z(n230) );
  CNIVX1 U237 ( .A(n232), .Z(n231) );
  CNIVX1 U238 ( .A(f02[11]), .Z(n232) );
  CNIVX1 U239 ( .A(n234), .Z(n233) );
  CNIVX1 U240 ( .A(n235), .Z(n234) );
  CNIVX1 U241 ( .A(f02[3]), .Z(n235) );
  CNIVX1 U242 ( .A(n237), .Z(n236) );
  CNIVX1 U243 ( .A(n238), .Z(n237) );
  CNIVX1 U244 ( .A(f02[7]), .Z(n238) );
  CNIVX1 U245 ( .A(n240), .Z(n239) );
  CNIVX1 U246 ( .A(n241), .Z(n240) );
  CNIVX1 U247 ( .A(f02[9]), .Z(n241) );
  CNIVX1 U248 ( .A(n243), .Z(n242) );
  CNIVX1 U249 ( .A(f02[19]), .Z(n243) );
  CNIVX1 U250 ( .A(n245), .Z(n244) );
  CNIVX1 U251 ( .A(f02[15]), .Z(n245) );
  CNIVX1 U252 ( .A(n247), .Z(n246) );
  CNIVX1 U253 ( .A(f02[17]), .Z(n247) );
  CNIVX1 U254 ( .A(captA[20]), .Z(n248) );
  CNIVX1 U255 ( .A(n710), .Z(n249) );
  CNIVX1 U256 ( .A(n518), .Z(n250) );
  CNIVX1 U257 ( .A(n252), .Z(n251) );
  CNIVX1 U258 ( .A(n253), .Z(n252) );
  CNIVX1 U259 ( .A(f11[1]), .Z(n253) );
  CNIVX1 U260 ( .A(n255), .Z(n254) );
  CNIVX1 U261 ( .A(n256), .Z(n255) );
  CNIVX1 U262 ( .A(f11[2]), .Z(n256) );
  CNIVX1 U263 ( .A(n258), .Z(n257) );
  CNIVX1 U264 ( .A(n259), .Z(n258) );
  CNIVX1 U265 ( .A(f21[2]), .Z(n259) );
  CNIVX1 U266 ( .A(n261), .Z(n260) );
  CNIVX1 U267 ( .A(f11[4]), .Z(n261) );
  CNIVX1 U268 ( .A(n263), .Z(n262) );
  CNIVX1 U269 ( .A(n264), .Z(n263) );
  CNIVX1 U270 ( .A(f11[3]), .Z(n264) );
  CNIVX1 U271 ( .A(n266), .Z(n265) );
  CNIVX1 U272 ( .A(f21[7]), .Z(n266) );
  CIVDX1 U273 ( .A(all_in1), .Z1(n268) );
  CNIVX1 U274 ( .A(n268), .Z(n267) );
  CIVDX1 U275 ( .A(all_in), .Z1(n270) );
  CNIVX1 U276 ( .A(n270), .Z(n269) );
  CNIVX1 U277 ( .A(n272), .Z(n271) );
  CNIVX1 U278 ( .A(captB[2]), .Z(n272) );
  CNIVX1 U279 ( .A(captB[23]), .Z(n273) );
  CNIVX1 U280 ( .A(n275), .Z(n274) );
  CNIVX1 U281 ( .A(n276), .Z(n275) );
  CNIVX1 U282 ( .A(n277), .Z(n276) );
  CNIVX1 U283 ( .A(f11[6]), .Z(n277) );
  CIVXL U284 ( .A(captA[17]), .Z(n278) );
  CIVX2 U285 ( .A(n278), .Z(n279) );
  CNIVX1 U286 ( .A(n281), .Z(n280) );
  CNIVX1 U287 ( .A(f21[13]), .Z(n281) );
  CNIVX1 U288 ( .A(n283), .Z(n282) );
  CNIVX1 U289 ( .A(f21[12]), .Z(n283) );
  CNIVX1 U290 ( .A(f01[4]), .Z(n284) );
  CIVDX1 U291 ( .A(all_in5), .Z1(n286) );
  CNIVX1 U292 ( .A(n286), .Z(n285) );
  CIVDX1 U293 ( .A(f15[27]), .Z1(n288) );
  CNIVX1 U294 ( .A(n288), .Z(n287) );
  CIVDX1 U295 ( .A(f15[22]), .Z1(n290) );
  CNIVX1 U296 ( .A(n290), .Z(n289) );
  CIVDX1 U297 ( .A(f15[17]), .Z1(n292) );
  CNIVX1 U298 ( .A(n292), .Z(n291) );
  CIVDX1 U299 ( .A(f15[12]), .Z1(n294) );
  CNIVX1 U300 ( .A(n294), .Z(n293) );
  CIVDX1 U301 ( .A(f15[7]), .Z1(n296) );
  CNIVX1 U302 ( .A(n296), .Z(n295) );
  CIVDX1 U303 ( .A(f15[2]), .Z1(n298) );
  CNIVX1 U304 ( .A(n298), .Z(n297) );
  CIVDX1 U305 ( .A(f23[30]), .Z1(n300) );
  CNIVX1 U306 ( .A(n300), .Z(n299) );
  CIVDX1 U307 ( .A(f23[25]), .Z1(n302) );
  CNIVX1 U308 ( .A(n302), .Z(n301) );
  CIVDX1 U309 ( .A(f23[20]), .Z1(n304) );
  CNIVX1 U310 ( .A(n304), .Z(n303) );
  CIVDX1 U311 ( .A(f23[15]), .Z1(n306) );
  CNIVX1 U312 ( .A(n306), .Z(n305) );
  CNIVX1 U313 ( .A(n1413), .Z(n307) );
  CNIVX1 U314 ( .A(n1408), .Z(n308) );
  CNIVX1 U315 ( .A(n1403), .Z(n309) );
  CNIVX1 U316 ( .A(n1398), .Z(n310) );
  CNIVX1 U317 ( .A(n1393), .Z(n311) );
  CNIVX1 U318 ( .A(n1388), .Z(n312) );
  CNIVX1 U319 ( .A(captB[26]), .Z(n313) );
  CNIVX1 U320 ( .A(n711), .Z(n314) );
  CNIVX1 U321 ( .A(n316), .Z(n315) );
  CNIVX1 U322 ( .A(n317), .Z(n316) );
  CNIVX1 U323 ( .A(f01[3]), .Z(n317) );
  CNIVX1 U324 ( .A(n363), .Z(n318) );
  CNIVX1 U325 ( .A(n320), .Z(n319) );
  CNIVX1 U326 ( .A(n650), .Z(n320) );
  CNIVX1 U327 ( .A(n322), .Z(n321) );
  CNIVX1 U328 ( .A(n323), .Z(n322) );
  CNIVX1 U329 ( .A(f01[7]), .Z(n323) );
  CNIVX1 U330 ( .A(n325), .Z(n324) );
  CNIVX1 U331 ( .A(captA[14]), .Z(n325) );
  CNIVX1 U332 ( .A(n202), .Z(n326) );
  CNIVX1 U333 ( .A(n328), .Z(n327) );
  CNIVX1 U334 ( .A(n329), .Z(n328) );
  CNIVX1 U335 ( .A(f21[3]), .Z(n329) );
  CNIVX1 U336 ( .A(n331), .Z(n330) );
  CNIVX1 U337 ( .A(n332), .Z(n331) );
  CNIVX1 U338 ( .A(captC[17]), .Z(n332) );
  CNIVX1 U339 ( .A(n334), .Z(n333) );
  CNIVX1 U340 ( .A(f01[17]), .Z(n334) );
  CNIVX1 U341 ( .A(n517), .Z(n335) );
  CIVDX1 U342 ( .A(f23[16]), .Z1(n337) );
  CNIVX1 U343 ( .A(n337), .Z(n336) );
  CIVDX1 U344 ( .A(f23[11]), .Z1(n339) );
  CNIVX1 U345 ( .A(n339), .Z(n338) );
  CIVDX1 U346 ( .A(f23[6]), .Z1(n341) );
  CNIVX1 U347 ( .A(n341), .Z(n340) );
  CIVDX1 U348 ( .A(f23[0]), .Z1(n343) );
  CNIVX1 U349 ( .A(n343), .Z(n342) );
  CIVDX1 U350 ( .A(f42[30]), .Z1(n345) );
  CNIVX1 U351 ( .A(n345), .Z(n344) );
  CIVDX1 U352 ( .A(f42[25]), .Z1(n347) );
  CNIVX1 U353 ( .A(n347), .Z(n346) );
  CIVDX1 U354 ( .A(f42[20]), .Z1(n349) );
  CNIVX1 U355 ( .A(n349), .Z(n348) );
  CIVDX1 U356 ( .A(f42[15]), .Z1(n351) );
  CNIVX1 U357 ( .A(n351), .Z(n350) );
  CIVDX1 U358 ( .A(f42[10]), .Z1(n353) );
  CNIVX1 U359 ( .A(n353), .Z(n352) );
  CIVDX1 U360 ( .A(f42[5]), .Z1(n355) );
  CNIVX1 U361 ( .A(n355), .Z(n354) );
  CIVDX1 U362 ( .A(f42[0]), .Z1(n357) );
  CNIVX1 U363 ( .A(n357), .Z(n356) );
  CNIVX1 U364 ( .A(n359), .Z(n358) );
  CNIVX1 U365 ( .A(n360), .Z(n359) );
  CNIVX1 U366 ( .A(f21[5]), .Z(n360) );
  CNIVX1 U367 ( .A(captA[23]), .Z(n361) );
  CNIVX1 U368 ( .A(captC[9]), .Z(n362) );
  CNIVX1 U369 ( .A(captB[9]), .Z(n363) );
  CIVDX1 U370 ( .A(f42[2]), .Z1(n365) );
  CNIVX1 U371 ( .A(n365), .Z(n364) );
  CIVDX1 U372 ( .A(f42[1]), .Z1(n367) );
  CNIVX1 U373 ( .A(n367), .Z(n366) );
  CIVDX1 U374 ( .A(f42[7]), .Z1(n369) );
  CNIVX1 U375 ( .A(n369), .Z(n368) );
  CIVDX1 U376 ( .A(f42[6]), .Z1(n371) );
  CNIVX1 U377 ( .A(n371), .Z(n370) );
  CIVDX1 U378 ( .A(f42[4]), .Z1(n373) );
  CNIVX1 U379 ( .A(n373), .Z(n372) );
  CIVDX1 U380 ( .A(f42[3]), .Z1(n375) );
  CNIVX1 U381 ( .A(n375), .Z(n374) );
  CIVDX1 U382 ( .A(f42[12]), .Z1(n377) );
  CNIVX1 U383 ( .A(n377), .Z(n376) );
  CIVDX1 U384 ( .A(f42[11]), .Z1(n379) );
  CNIVX1 U385 ( .A(n379), .Z(n378) );
  CIVDX1 U386 ( .A(f42[9]), .Z1(n381) );
  CNIVX1 U387 ( .A(n381), .Z(n380) );
  CIVDX1 U388 ( .A(f42[8]), .Z1(n383) );
  CNIVX1 U389 ( .A(n383), .Z(n382) );
  CIVDX1 U390 ( .A(f42[17]), .Z1(n385) );
  CNIVX1 U391 ( .A(n385), .Z(n384) );
  CIVDX1 U392 ( .A(f42[16]), .Z1(n387) );
  CNIVX1 U393 ( .A(n387), .Z(n386) );
  CIVDX1 U394 ( .A(f42[14]), .Z1(n389) );
  CNIVX1 U395 ( .A(n389), .Z(n388) );
  CIVDX1 U396 ( .A(f42[13]), .Z1(n391) );
  CNIVX1 U397 ( .A(n391), .Z(n390) );
  CIVDX1 U398 ( .A(f42[22]), .Z1(n393) );
  CNIVX1 U399 ( .A(n393), .Z(n392) );
  CIVDX1 U400 ( .A(f42[21]), .Z1(n395) );
  CNIVX1 U401 ( .A(n395), .Z(n394) );
  CIVDX1 U402 ( .A(f42[19]), .Z1(n397) );
  CNIVX1 U403 ( .A(n397), .Z(n396) );
  CIVDX1 U404 ( .A(f42[18]), .Z1(n399) );
  CNIVX1 U405 ( .A(n399), .Z(n398) );
  CIVDX1 U406 ( .A(f42[27]), .Z1(n401) );
  CNIVX1 U407 ( .A(n401), .Z(n400) );
  CIVDX1 U408 ( .A(f42[26]), .Z1(n403) );
  CNIVX1 U409 ( .A(n403), .Z(n402) );
  CIVDX1 U410 ( .A(f42[24]), .Z1(n405) );
  CNIVX1 U411 ( .A(n405), .Z(n404) );
  CIVDX1 U412 ( .A(f42[23]), .Z1(n407) );
  CNIVX1 U413 ( .A(n407), .Z(n406) );
  CIVDX1 U414 ( .A(f42[31]), .Z1(n409) );
  CNIVX1 U415 ( .A(n409), .Z(n408) );
  CIVDX1 U416 ( .A(f42[29]), .Z1(n411) );
  CNIVX1 U417 ( .A(n411), .Z(n410) );
  CIVDX1 U418 ( .A(f42[28]), .Z1(n413) );
  CNIVX1 U419 ( .A(n413), .Z(n412) );
  CIVDX1 U420 ( .A(f23[3]), .Z1(n415) );
  CNIVX1 U421 ( .A(n415), .Z(n414) );
  CIVDX1 U422 ( .A(f23[2]), .Z1(n417) );
  CNIVX1 U423 ( .A(n417), .Z(n416) );
  CIVDX1 U424 ( .A(f23[8]), .Z1(n419) );
  CNIVX1 U425 ( .A(n419), .Z(n418) );
  CIVDX1 U426 ( .A(f23[7]), .Z1(n421) );
  CNIVX1 U427 ( .A(n421), .Z(n420) );
  CIVDX1 U428 ( .A(f23[5]), .Z1(n423) );
  CNIVX1 U429 ( .A(n423), .Z(n422) );
  CIVDX1 U430 ( .A(f23[4]), .Z1(n425) );
  CNIVX1 U431 ( .A(n425), .Z(n424) );
  CIVDX1 U432 ( .A(f23[13]), .Z1(n427) );
  CNIVX1 U433 ( .A(n427), .Z(n426) );
  CIVDX1 U434 ( .A(f23[12]), .Z1(n429) );
  CNIVX1 U435 ( .A(n429), .Z(n428) );
  CIVDX1 U436 ( .A(f23[10]), .Z1(n431) );
  CNIVX1 U437 ( .A(n431), .Z(n430) );
  CIVDX1 U438 ( .A(f23[9]), .Z1(n433) );
  CNIVX1 U439 ( .A(n433), .Z(n432) );
  CIVDX1 U440 ( .A(f23[18]), .Z1(n435) );
  CNIVX1 U441 ( .A(n435), .Z(n434) );
  CIVDX1 U442 ( .A(f23[17]), .Z1(n437) );
  CNIVX1 U443 ( .A(n437), .Z(n436) );
  CNIVX1 U444 ( .A(n439), .Z(n438) );
  CNIVX1 U445 ( .A(n440), .Z(n439) );
  CNIVX1 U446 ( .A(f01[21]), .Z(n440) );
  CNIVX1 U447 ( .A(captA[21]), .Z(n441) );
  CNIVX1 U448 ( .A(n443), .Z(n442) );
  CNIVX1 U449 ( .A(captA[2]), .Z(n443) );
  CNIVX1 U450 ( .A(f01[12]), .Z(n444) );
  CNIVX1 U451 ( .A(n446), .Z(n445) );
  CNIVX1 U452 ( .A(f02[6]), .Z(n446) );
  CNIVX1 U453 ( .A(n448), .Z(n447) );
  CNIVX1 U454 ( .A(captB[6]), .Z(n448) );
  CNIVX1 U455 ( .A(n450), .Z(n449) );
  CNIVX1 U456 ( .A(n451), .Z(n450) );
  CNIVX1 U457 ( .A(f21[4]), .Z(n451) );
  CNIVX1 U458 ( .A(n453), .Z(n452) );
  CNIVX1 U459 ( .A(captA[9]), .Z(n453) );
  CNIVX1 U460 ( .A(n455), .Z(n454) );
  CNIVX1 U461 ( .A(captA[8]), .Z(n455) );
  CNIVX1 U462 ( .A(f01[6]), .Z(n456) );
  CNIVX1 U463 ( .A(n458), .Z(n457) );
  CNIVX1 U464 ( .A(captA[6]), .Z(n458) );
  CNIVX1 U465 ( .A(captB[21]), .Z(n459) );
  CNIVX1 U466 ( .A(n461), .Z(n460) );
  CNIVX1 U467 ( .A(n462), .Z(n461) );
  CNIVX1 U468 ( .A(f02[1]), .Z(n462) );
  CNIVX1 U469 ( .A(n516), .Z(n463) );
  CNIVX1 U470 ( .A(n465), .Z(n464) );
  CNIVX1 U471 ( .A(n514), .Z(n465) );
  CNIVX1 U472 ( .A(n467), .Z(n466) );
  CNIVX1 U473 ( .A(f11[5]), .Z(n467) );
  CNIVX1 U474 ( .A(n469), .Z(n468) );
  CNIVX1 U475 ( .A(n470), .Z(n469) );
  CNIVX1 U476 ( .A(f11[0]), .Z(n470) );
  CNIVX1 U477 ( .A(n472), .Z(n471) );
  CNIVX1 U478 ( .A(f01[0]), .Z(n472) );
  CNIVX1 U479 ( .A(n474), .Z(n473) );
  CNIVX1 U480 ( .A(n475), .Z(n474) );
  CNIVX1 U481 ( .A(f21[1]), .Z(n475) );
  CNIVX1 U482 ( .A(n477), .Z(n476) );
  CNIVX1 U483 ( .A(n478), .Z(n477) );
  CNIVX1 U484 ( .A(f02[23]), .Z(n478) );
  CNIVX1 U485 ( .A(f01[2]), .Z(n479) );
  CNIVX1 U486 ( .A(n481), .Z(n480) );
  CNIVX1 U487 ( .A(captC[2]), .Z(n481) );
  CNIVX1 U488 ( .A(n712), .Z(n482) );
  CIVX2 U489 ( .A(n503), .Z(n483) );
  CIVX2 U490 ( .A(n483), .Z(n484) );
  CNIVX1 U491 ( .A(n486), .Z(n485) );
  CNIVX1 U492 ( .A(captA[7]), .Z(n486) );
  CNIVX1 U493 ( .A(n488), .Z(n487) );
  CNIVX1 U494 ( .A(captB[7]), .Z(n488) );
  CNIVX1 U495 ( .A(n490), .Z(n489) );
  CNIVX1 U496 ( .A(f02[8]), .Z(n490) );
  CNIVX1 U497 ( .A(n492), .Z(n491) );
  CNIVX1 U498 ( .A(captB[8]), .Z(n492) );
  CNIVX1 U499 ( .A(n494), .Z(n493) );
  CNIVX1 U500 ( .A(n495), .Z(n494) );
  CNIVX1 U501 ( .A(f01[19]), .Z(n495) );
  CNIVX1 U502 ( .A(n497), .Z(n496) );
  CNIVX1 U503 ( .A(n498), .Z(n497) );
  CNIVX1 U504 ( .A(captA[19]), .Z(n498) );
  CNIVX1 U505 ( .A(n500), .Z(n499) );
  CNIVX1 U506 ( .A(captA[5]), .Z(n500) );
  CNIVX1 U507 ( .A(n521), .Z(n501) );
  CIVX2 U508 ( .A(n504), .Z(n502) );
  CNIVX1 U509 ( .A(captA[0]), .Z(n504) );
  CNIVX1 U510 ( .A(n506), .Z(n505) );
  CNIVX1 U511 ( .A(n519), .Z(n506) );
  CNIVX1 U512 ( .A(n508), .Z(n507) );
  CNIVX1 U513 ( .A(n520), .Z(n508) );
  CNIVX1 U514 ( .A(n510), .Z(n509) );
  CNIVX1 U515 ( .A(n511), .Z(n510) );
  CNIVX1 U516 ( .A(captC[11]), .Z(n511) );
  CNIVX1 U517 ( .A(captC[23]), .Z(n512) );
  CNIVX1 U518 ( .A(captB[24]), .Z(n513) );
  CNIVX1 U519 ( .A(captB[14]), .Z(n514) );
  CNIVX1 U520 ( .A(captB[3]), .Z(n515) );
  CNIVX1 U521 ( .A(captB[11]), .Z(n516) );
  CNIVX1 U522 ( .A(captA[12]), .Z(n517) );
  CNIVX1 U523 ( .A(captA[11]), .Z(n518) );
  CNIVX1 U524 ( .A(captA[15]), .Z(n519) );
  CNIVX1 U525 ( .A(captA[13]), .Z(n520) );
  CNIVX1 U526 ( .A(captB[13]), .Z(n521) );
  CNIVX1 U527 ( .A(n523), .Z(n522) );
  CNIVX1 U528 ( .A(captA[4]), .Z(n523) );
  CNIVX1 U529 ( .A(n527), .Z(n524) );
  CIVX2 U530 ( .A(captC[0]), .Z(n525) );
  CIVX2 U531 ( .A(n525), .Z(n526) );
  CNIVX1 U532 ( .A(n529), .Z(n528) );
  CNIVX1 U533 ( .A(n530), .Z(n529) );
  CNIVX1 U534 ( .A(captA[16]), .Z(n530) );
  CNIVX1 U535 ( .A(n532), .Z(n531) );
  CNIVX1 U536 ( .A(n533), .Z(n532) );
  CNIVX1 U537 ( .A(captA[10]), .Z(n533) );
  CNIVX1 U538 ( .A(n535), .Z(n534) );
  CNIVX1 U539 ( .A(f11[10]), .Z(n535) );
  CNIVX1 U540 ( .A(n537), .Z(n536) );
  CNIVX1 U541 ( .A(f11[9]), .Z(n537) );
  CNIVX1 U542 ( .A(n1390), .Z(n538) );
  CNIVX1 U543 ( .A(n1384), .Z(n539) );
  CNIVX1 U544 ( .A(n1385), .Z(n540) );
  CNIVX1 U545 ( .A(n1395), .Z(n541) );
  CNIVX1 U546 ( .A(n1386), .Z(n542) );
  CNIVX1 U547 ( .A(n1387), .Z(n543) );
  CNIVX1 U548 ( .A(n1389), .Z(n544) );
  CNIVX1 U549 ( .A(n1400), .Z(n545) );
  CNIVX1 U550 ( .A(n1391), .Z(n546) );
  CNIVX1 U551 ( .A(n1392), .Z(n547) );
  CNIVX1 U552 ( .A(n1394), .Z(n548) );
  CNIVX1 U553 ( .A(n1405), .Z(n549) );
  CNIVX1 U554 ( .A(n1396), .Z(n550) );
  CNIVX1 U555 ( .A(n1397), .Z(n551) );
  CNIVX1 U556 ( .A(n1399), .Z(n552) );
  CNIVX1 U557 ( .A(n1410), .Z(n553) );
  CNIVX1 U558 ( .A(n1401), .Z(n554) );
  CNIVX1 U559 ( .A(n1402), .Z(n555) );
  CNIVX1 U560 ( .A(n1404), .Z(n556) );
  CNIVX1 U561 ( .A(n1415), .Z(n557) );
  CNIVX1 U562 ( .A(n1406), .Z(n558) );
  CNIVX1 U563 ( .A(n1407), .Z(n559) );
  CNIVX1 U564 ( .A(n1409), .Z(n560) );
  CIVDX1 U565 ( .A(all_in9), .Z1(n562) );
  CNIVX1 U566 ( .A(n562), .Z(n561) );
  CNIVX1 U567 ( .A(n1411), .Z(n563) );
  CNIVX1 U568 ( .A(n1412), .Z(n564) );
  CNIVX1 U569 ( .A(n1414), .Z(n565) );
  CIVDX1 U570 ( .A(f23[14]), .Z1(n567) );
  CNIVX1 U571 ( .A(n567), .Z(n566) );
  CIVDX1 U572 ( .A(f23[23]), .Z1(n569) );
  CNIVX1 U573 ( .A(n569), .Z(n568) );
  CIVDX1 U574 ( .A(f23[22]), .Z1(n571) );
  CNIVX1 U575 ( .A(n571), .Z(n570) );
  CIVDX1 U576 ( .A(f23[21]), .Z1(n573) );
  CNIVX1 U577 ( .A(n573), .Z(n572) );
  CIVDX1 U578 ( .A(f23[19]), .Z1(n575) );
  CNIVX1 U579 ( .A(n575), .Z(n574) );
  CIVDX1 U580 ( .A(f23[28]), .Z1(n577) );
  CNIVX1 U581 ( .A(n577), .Z(n576) );
  CIVDX1 U582 ( .A(f23[27]), .Z1(n579) );
  CNIVX1 U583 ( .A(n579), .Z(n578) );
  CIVDX1 U584 ( .A(f23[26]), .Z1(n581) );
  CNIVX1 U585 ( .A(n581), .Z(n580) );
  CIVDX1 U586 ( .A(f23[24]), .Z1(n583) );
  CNIVX1 U587 ( .A(n583), .Z(n582) );
  CIVDX1 U588 ( .A(f23[31]), .Z1(n585) );
  CNIVX1 U589 ( .A(n585), .Z(n584) );
  CIVDX1 U590 ( .A(f23[29]), .Z1(n587) );
  CNIVX1 U591 ( .A(n587), .Z(n586) );
  CIVDX1 U592 ( .A(f15[5]), .Z1(n589) );
  CNIVX1 U593 ( .A(n589), .Z(n588) );
  CIVDX1 U594 ( .A(f15[4]), .Z1(n591) );
  CNIVX1 U595 ( .A(n591), .Z(n590) );
  CIVDX1 U596 ( .A(f15[3]), .Z1(n593) );
  CNIVX1 U597 ( .A(n593), .Z(n592) );
  CIVDX1 U598 ( .A(f15[0]), .Z1(n595) );
  CNIVX1 U599 ( .A(n595), .Z(n594) );
  CIVDX1 U600 ( .A(f15[10]), .Z1(n597) );
  CNIVX1 U601 ( .A(n597), .Z(n596) );
  CIVDX1 U602 ( .A(f15[9]), .Z1(n599) );
  CNIVX1 U603 ( .A(n599), .Z(n598) );
  CIVDX1 U604 ( .A(f15[8]), .Z1(n601) );
  CNIVX1 U605 ( .A(n601), .Z(n600) );
  CIVDX1 U606 ( .A(f15[6]), .Z1(n603) );
  CNIVX1 U607 ( .A(n603), .Z(n602) );
  CIVDX1 U608 ( .A(f15[15]), .Z1(n605) );
  CNIVX1 U609 ( .A(n605), .Z(n604) );
  CIVDX1 U610 ( .A(f15[14]), .Z1(n607) );
  CNIVX1 U611 ( .A(n607), .Z(n606) );
  CIVDX1 U612 ( .A(f15[13]), .Z1(n609) );
  CNIVX1 U613 ( .A(n609), .Z(n608) );
  CIVDX1 U614 ( .A(f15[11]), .Z1(n611) );
  CNIVX1 U615 ( .A(n611), .Z(n610) );
  CIVDX1 U616 ( .A(f15[20]), .Z1(n613) );
  CNIVX1 U617 ( .A(n613), .Z(n612) );
  CIVDX1 U618 ( .A(f15[19]), .Z1(n615) );
  CNIVX1 U619 ( .A(n615), .Z(n614) );
  CIVDX1 U620 ( .A(f15[18]), .Z1(n617) );
  CNIVX1 U621 ( .A(n617), .Z(n616) );
  CIVDX1 U622 ( .A(f15[16]), .Z1(n619) );
  CNIVX1 U623 ( .A(n619), .Z(n618) );
  CIVDX1 U624 ( .A(f15[25]), .Z1(n621) );
  CNIVX1 U625 ( .A(n621), .Z(n620) );
  CIVDX1 U626 ( .A(f15[24]), .Z1(n623) );
  CNIVX1 U627 ( .A(n623), .Z(n622) );
  CIVDX1 U628 ( .A(f15[23]), .Z1(n625) );
  CNIVX1 U629 ( .A(n625), .Z(n624) );
  CIVDX1 U630 ( .A(f15[21]), .Z1(n627) );
  CNIVX1 U631 ( .A(n627), .Z(n626) );
  CIVDX1 U632 ( .A(f15[30]), .Z1(n629) );
  CNIVX1 U633 ( .A(n629), .Z(n628) );
  CIVDX1 U634 ( .A(f15[29]), .Z1(n631) );
  CNIVX1 U635 ( .A(n631), .Z(n630) );
  CIVDX1 U636 ( .A(f15[28]), .Z1(n633) );
  CNIVX1 U637 ( .A(n633), .Z(n632) );
  CIVDX1 U638 ( .A(f15[26]), .Z1(n635) );
  CNIVX1 U639 ( .A(n635), .Z(n634) );
  CIVDX1 U640 ( .A(f15[31]), .Z1(n637) );
  CNIVX1 U641 ( .A(n637), .Z(n636) );
  CIVDX1 U642 ( .A(all_in7), .Z1(n639) );
  CNIVX1 U643 ( .A(n639), .Z(n638) );
  CIVDX1 U644 ( .A(all_in8), .Z1(n641) );
  CNIVX1 U645 ( .A(n641), .Z(n640) );
  CIVDX1 U646 ( .A(all_in2), .Z1(n643) );
  CNIVX1 U647 ( .A(n643), .Z(n642) );
  CIVDX1 U648 ( .A(all_in3), .Z1(n645) );
  CNIVX1 U649 ( .A(n645), .Z(n644) );
  CIVDX1 U650 ( .A(all_in4), .Z1(n647) );
  CNIVX1 U651 ( .A(n647), .Z(n646) );
  CIVDX1 U652 ( .A(all_in6), .Z1(n649) );
  CNIVX1 U653 ( .A(n649), .Z(n648) );
  CNIVX1 U654 ( .A(captC[14]), .Z(n650) );
  CNIVX1 U655 ( .A(n652), .Z(n651) );
  CNIVX1 U656 ( .A(captC[3]), .Z(n652) );
  CNIVX1 U657 ( .A(n654), .Z(n653) );
  CNIVX1 U658 ( .A(captC[4]), .Z(n654) );
  CNIVX1 U659 ( .A(n656), .Z(n655) );
  CNIVX1 U660 ( .A(captC[5]), .Z(n656) );
  CNIVX1 U661 ( .A(n658), .Z(n657) );
  CNIVX1 U662 ( .A(captC[12]), .Z(n658) );
  CNIVX1 U663 ( .A(n660), .Z(n659) );
  CNIVX1 U664 ( .A(n661), .Z(n660) );
  CNIVX1 U665 ( .A(captC[13]), .Z(n661) );
  CNIVX1 U666 ( .A(n663), .Z(n662) );
  CNIVX1 U667 ( .A(n664), .Z(n663) );
  CNIVX1 U668 ( .A(captC[15]), .Z(n664) );
  CNIVX1 U669 ( .A(n666), .Z(n665) );
  CNIVX1 U670 ( .A(n667), .Z(n666) );
  CNIVX1 U671 ( .A(captC[16]), .Z(n667) );
  CNIVX1 U672 ( .A(n669), .Z(n668) );
  CNIVX1 U673 ( .A(n670), .Z(n669) );
  CNIVX1 U674 ( .A(captC[18]), .Z(n670) );
  CNIVX1 U675 ( .A(n672), .Z(n671) );
  CNIVX1 U676 ( .A(n673), .Z(n672) );
  CNIVX1 U677 ( .A(captC[19]), .Z(n673) );
  CNIVX1 U678 ( .A(n675), .Z(n674) );
  CNIVX1 U679 ( .A(n676), .Z(n675) );
  CNIVX1 U680 ( .A(captC[20]), .Z(n676) );
  CNIVX1 U681 ( .A(captC[21]), .Z(n677) );
  CNIVX1 U682 ( .A(n680), .Z(n678) );
  CIVX2 U683 ( .A(n681), .Z(n679) );
  CIVX2 U684 ( .A(n679), .Z(n680) );
  CNIVX1 U685 ( .A(captB[0]), .Z(n681) );
  CNIVX1 U686 ( .A(n683), .Z(n682) );
  CNIVX1 U687 ( .A(captB[5]), .Z(n683) );
  CNIVX1 U688 ( .A(n685), .Z(n684) );
  CNIVX1 U689 ( .A(captB[10]), .Z(n685) );
  CNIVX1 U690 ( .A(n687), .Z(n686) );
  CNIVX1 U691 ( .A(captB[12]), .Z(n687) );
  CNIVX1 U692 ( .A(n689), .Z(n688) );
  CNIVX1 U693 ( .A(n690), .Z(n689) );
  CNIVX1 U694 ( .A(captB[15]), .Z(n690) );
  CNIVX1 U695 ( .A(n692), .Z(n691) );
  CNIVX1 U696 ( .A(n693), .Z(n692) );
  CNIVX1 U697 ( .A(captB[16]), .Z(n693) );
  CNIVX1 U698 ( .A(n695), .Z(n694) );
  CNIVX1 U699 ( .A(n696), .Z(n695) );
  CNIVX1 U700 ( .A(captB[18]), .Z(n696) );
  CNIVX1 U701 ( .A(n698), .Z(n697) );
  CNIVX1 U702 ( .A(n699), .Z(n698) );
  CNIVX1 U703 ( .A(captB[19]), .Z(n699) );
  CNIVX1 U704 ( .A(n701), .Z(n700) );
  CNIVX1 U705 ( .A(n702), .Z(n701) );
  CNIVX1 U706 ( .A(captB[20]), .Z(n702) );
  CNIVX1 U707 ( .A(captB[22]), .Z(n703) );
  CNIVX1 U708 ( .A(captB[25]), .Z(n704) );
  CNIVX1 U709 ( .A(captB[27]), .Z(n705) );
  CNIVX1 U710 ( .A(captB[29]), .Z(n706) );
  CNIVX1 U711 ( .A(n708), .Z(n707) );
  CNIVX1 U712 ( .A(captA[3]), .Z(n708) );
  CNIVX1 U713 ( .A(captA[27]), .Z(n709) );
  CNIVX1 U714 ( .A(captC[1]), .Z(n710) );
  CNIVX1 U715 ( .A(captB[1]), .Z(n711) );
  CNIVX1 U716 ( .A(captA[1]), .Z(n712) );
  CNIVX1 U717 ( .A(n714), .Z(n713) );
  CNIVX1 U718 ( .A(f02[18]), .Z(n714) );
  CNIVX1 U719 ( .A(n716), .Z(n715) );
  CNIVX1 U720 ( .A(f02[16]), .Z(n716) );
  CNIVXL U721 ( .A(captA[31]), .Z(n1378) );
  CNIVX1 U722 ( .A(n1378), .Z(n717) );
  CNIVX1 U723 ( .A(n719), .Z(n718) );
  CNIVX1 U724 ( .A(f02[20]), .Z(n719) );
  CNIVX1 U725 ( .A(n721), .Z(n720) );
  CNIVX1 U726 ( .A(captC[10]), .Z(n721) );
  CNIVX1 U727 ( .A(n723), .Z(n722) );
  CNIVX1 U728 ( .A(captC[27]), .Z(n723) );
  CNIVXL U729 ( .A(captB[31]), .Z(n1379) );
  CNIVX1 U730 ( .A(n1379), .Z(n724) );
  CNIVX1 U731 ( .A(n726), .Z(n725) );
  CNIVX1 U732 ( .A(f02[22]), .Z(n726) );
  CNIVX1 U733 ( .A(n728), .Z(n727) );
  CNIVX1 U734 ( .A(captC[26]), .Z(n728) );
  CNIVX1 U735 ( .A(n730), .Z(n729) );
  CNIVX1 U736 ( .A(captA[24]), .Z(n730) );
  CNIVX1 U737 ( .A(n732), .Z(n731) );
  CNIVX1 U738 ( .A(captA[22]), .Z(n732) );
  CNIVX1 U739 ( .A(n734), .Z(n733) );
  CNIVX1 U740 ( .A(n735), .Z(n734) );
  CNIVX1 U741 ( .A(captA[18]), .Z(n735) );
  CNIVX1 U742 ( .A(n737), .Z(n736) );
  CNIVX1 U743 ( .A(captB[28]), .Z(n737) );
  CIVDX1 U744 ( .A(captA[30]), .Z1(n738) );
  CNIVX1 U745 ( .A(n740), .Z(n739) );
  CNIVX1 U746 ( .A(captA[28]), .Z(n740) );
  CNIVX1 U747 ( .A(n742), .Z(n741) );
  CNIVX1 U748 ( .A(captA[26]), .Z(n742) );
  CNIVX1 U749 ( .A(n744), .Z(n743) );
  CNIVX1 U750 ( .A(f02[25]), .Z(n744) );
  CNIVX1 U751 ( .A(n746), .Z(n745) );
  CNIVX1 U752 ( .A(f02[24]), .Z(n746) );
  CNIVX1 U753 ( .A(n748), .Z(n747) );
  CNIVX1 U754 ( .A(f11[21]), .Z(n748) );
  CNIVX1 U755 ( .A(n750), .Z(n749) );
  CNIVX1 U756 ( .A(f11[16]), .Z(n750) );
  CNIVX1 U757 ( .A(n752), .Z(n751) );
  CNIVX1 U758 ( .A(n753), .Z(n752) );
  CNIVX1 U759 ( .A(f11[22]), .Z(n753) );
  CNIVX1 U760 ( .A(n755), .Z(n754) );
  CNIVX1 U761 ( .A(f11[18]), .Z(n755) );
  CNIVX1 U762 ( .A(n757), .Z(n756) );
  CNIVX1 U763 ( .A(captC[29]), .Z(n757) );
  CNIVX1 U764 ( .A(n759), .Z(n758) );
  CNIVX1 U765 ( .A(captC[28]), .Z(n759) );
  CIVDX1 U766 ( .A(captB[30]), .Z1(n760) );
  CNIVX1 U767 ( .A(n762), .Z(n761) );
  CNIVX1 U768 ( .A(n763), .Z(n762) );
  CNIVX1 U769 ( .A(f01[23]), .Z(n763) );
  CNIVX1 U770 ( .A(f02[27]), .Z(n764) );
  CNIVX1 U771 ( .A(n766), .Z(n765) );
  CNIVX1 U772 ( .A(f02[26]), .Z(n766) );
  CNIVX1 U773 ( .A(n768), .Z(n767) );
  CNIVX1 U774 ( .A(f11[19]), .Z(n768) );
  CNIVX1 U775 ( .A(n770), .Z(n769) );
  CNIVX1 U776 ( .A(f01[25]), .Z(n770) );
  CNIVX1 U777 ( .A(n772), .Z(n771) );
  CNIVX1 U778 ( .A(f11[20]), .Z(n772) );
  CNIVX1 U779 ( .A(f01[24]), .Z(n773) );
  CNIVX1 U780 ( .A(n775), .Z(n774) );
  CNIVX1 U781 ( .A(f11[17]), .Z(n775) );
  CNIVX1 U782 ( .A(f11[27]), .Z(n776) );
  CNIVX1 U783 ( .A(f11[26]), .Z(n777) );
  CNIVX1 U784 ( .A(f21[27]), .Z(n778) );
  CIVDX1 U785 ( .A(captC[30]), .Z1(n779) );
  CNIVX1 U786 ( .A(n781), .Z(n780) );
  CNIVX1 U787 ( .A(f02[29]), .Z(n781) );
  CNIVX1 U788 ( .A(n784), .Z(n783) );
  CNIVX1 U789 ( .A(n785), .Z(n784) );
  CNIVX1 U790 ( .A(f02[0]), .Z(n785) );
  CNIVX1 U791 ( .A(f21[24]), .Z(n786) );
  CNIVX1 U792 ( .A(f01[27]), .Z(n787) );
  CNIVX1 U793 ( .A(f01[26]), .Z(n788) );
  CNIVX1 U794 ( .A(n790), .Z(n789) );
  CNIVX1 U795 ( .A(f11[29]), .Z(n790) );
  CNIVX1 U796 ( .A(n792), .Z(n791) );
  CNIVX1 U797 ( .A(f11[28]), .Z(n792) );
  CNIVX1 U798 ( .A(f21[26]), .Z(n793) );
  CDLY1XL U799 ( .A(f11[8]), .Z(n794) );
  CNIVX1 U800 ( .A(n796), .Z(n795) );
  CNIVX1 U801 ( .A(n797), .Z(n796) );
  CNIVX1 U802 ( .A(f11[7]), .Z(n797) );
  CNIVX1 U803 ( .A(n799), .Z(n798) );
  CNIVX1 U804 ( .A(n800), .Z(n799) );
  CNIVX1 U805 ( .A(n801), .Z(n800) );
  CNIVX1 U806 ( .A(f11[12]), .Z(n801) );
  CDLY1XL U807 ( .A(f11[11]), .Z(n802) );
  CNIVX1 U808 ( .A(n804), .Z(n803) );
  CNIVX1 U809 ( .A(n805), .Z(n804) );
  CNIVX1 U810 ( .A(f01[5]), .Z(n805) );
  CNIVX1 U811 ( .A(n807), .Z(n806) );
  CNIVX1 U812 ( .A(f01[15]), .Z(n807) );
  CNIVX1 U813 ( .A(n809), .Z(n808) );
  CNIVX1 U814 ( .A(f01[8]), .Z(n809) );
  CNIVX1 U815 ( .A(n811), .Z(n810) );
  CNIVX1 U816 ( .A(f01[13]), .Z(n811) );
  CDLY1XL U817 ( .A(f11[13]), .Z(n812) );
  CNIVX1 U818 ( .A(n814), .Z(n813) );
  CNIVX1 U819 ( .A(n815), .Z(n814) );
  CNIVX1 U820 ( .A(f01[11]), .Z(n815) );
  CNIVX1 U821 ( .A(n817), .Z(n816) );
  CNIVX1 U822 ( .A(n818), .Z(n817) );
  CNIVX1 U823 ( .A(f01[9]), .Z(n818) );
  CNIVX1 U824 ( .A(n820), .Z(n819) );
  CNIVX1 U825 ( .A(f11[15]), .Z(n820) );
  CNIVX1 U826 ( .A(n822), .Z(n821) );
  CNIVX1 U827 ( .A(n823), .Z(n822) );
  CNIVX1 U828 ( .A(n824), .Z(n823) );
  CNIVX1 U829 ( .A(f11[14]), .Z(n824) );
  CIVDX1 U830 ( .A(f37[9]), .Z1(n826) );
  CNIVX1 U831 ( .A(n826), .Z(n825) );
  CIVDX1 U832 ( .A(f54[9]), .Z1(n828) );
  CNIVX1 U833 ( .A(n828), .Z(n827) );
  CNIVXL U834 ( .A(captC[31]), .Z(n1380) );
  CNIVX1 U835 ( .A(n1380), .Z(n829) );
  CNIVX2 U836 ( .A(f21[28]), .Z(n830) );
  CIVDX1 U837 ( .A(f54[20]), .Z1(n832) );
  CNIVX1 U838 ( .A(n832), .Z(n831) );
  CIVDX1 U839 ( .A(f54[18]), .Z1(n834) );
  CNIVX1 U840 ( .A(n834), .Z(n833) );
  CIVDX1 U841 ( .A(f54[6]), .Z1(n836) );
  CNIVX1 U842 ( .A(n836), .Z(n835) );
  CIVDX1 U843 ( .A(f54[2]), .Z1(n838) );
  CNIVX1 U844 ( .A(n838), .Z(n837) );
  CIVDX1 U845 ( .A(f54[22]), .Z1(n840) );
  CNIVX1 U846 ( .A(n840), .Z(n839) );
  CIVDX1 U847 ( .A(f37[20]), .Z1(n842) );
  CNIVX1 U848 ( .A(n842), .Z(n841) );
  CIVDX1 U849 ( .A(f37[18]), .Z1(n844) );
  CNIVX1 U850 ( .A(n844), .Z(n843) );
  CIVDX1 U851 ( .A(f37[6]), .Z1(n846) );
  CNIVX1 U852 ( .A(n846), .Z(n845) );
  CIVDX1 U853 ( .A(f37[2]), .Z1(n848) );
  CNIVX1 U854 ( .A(n848), .Z(n847) );
  CIVDX1 U855 ( .A(f37[22]), .Z1(n850) );
  CNIVX1 U856 ( .A(n850), .Z(n849) );
  CIVDX1 U857 ( .A(f37[12]), .Z1(n852) );
  CNIVX1 U858 ( .A(n852), .Z(n851) );
  CIVDX1 U859 ( .A(f54[12]), .Z1(n854) );
  CNIVX1 U860 ( .A(n854), .Z(n853) );
  CIVDX1 U861 ( .A(f54[10]), .Z1(n856) );
  CNIVX1 U862 ( .A(n856), .Z(n855) );
  CIVDX1 U863 ( .A(f37[14]), .Z1(n858) );
  CNIVX1 U864 ( .A(n858), .Z(n857) );
  CIVDX1 U865 ( .A(f54[14]), .Z1(n860) );
  CNIVX1 U866 ( .A(n860), .Z(n859) );
  CIVDX1 U867 ( .A(f37[10]), .Z1(n862) );
  CNIVX1 U868 ( .A(n862), .Z(n861) );
  CIVDX1 U869 ( .A(f54[8]), .Z1(n864) );
  CNIVX1 U870 ( .A(n864), .Z(n863) );
  CIVDX1 U871 ( .A(f54[5]), .Z1(n866) );
  CNIVX1 U872 ( .A(n866), .Z(n865) );
  CIVDX1 U873 ( .A(f54[4]), .Z1(n868) );
  CNIVX1 U874 ( .A(n868), .Z(n867) );
  CIVDX1 U875 ( .A(f54[23]), .Z1(n870) );
  CNIVX1 U876 ( .A(n870), .Z(n869) );
  CIVDX1 U877 ( .A(f54[21]), .Z1(n872) );
  CNIVX1 U878 ( .A(n872), .Z(n871) );
  CIVDX1 U879 ( .A(f54[19]), .Z1(n874) );
  CNIVX1 U880 ( .A(n874), .Z(n873) );
  CIVDX1 U881 ( .A(f54[17]), .Z1(n876) );
  CNIVX1 U882 ( .A(n876), .Z(n875) );
  CIVDX1 U883 ( .A(f54[16]), .Z1(n878) );
  CNIVX1 U884 ( .A(n878), .Z(n877) );
  CIVDX1 U885 ( .A(f37[5]), .Z1(n880) );
  CNIVX1 U886 ( .A(n880), .Z(n879) );
  CIVDX1 U887 ( .A(f37[4]), .Z1(n882) );
  CNIVX1 U888 ( .A(n882), .Z(n881) );
  CIVDX1 U889 ( .A(f37[21]), .Z1(n884) );
  CNIVX1 U890 ( .A(n884), .Z(n883) );
  CIVDX1 U891 ( .A(f37[19]), .Z1(n886) );
  CNIVX1 U892 ( .A(n886), .Z(n885) );
  CIVDX1 U893 ( .A(f37[17]), .Z1(n888) );
  CNIVX1 U894 ( .A(n888), .Z(n887) );
  CIVDX1 U895 ( .A(f37[16]), .Z1(n890) );
  CNIVX1 U896 ( .A(n890), .Z(n889) );
  CIVDX1 U897 ( .A(f37[8]), .Z1(n892) );
  CNIVX1 U898 ( .A(n892), .Z(n891) );
  CIVDX1 U899 ( .A(f37[23]), .Z1(n894) );
  CNIVX1 U900 ( .A(n894), .Z(n893) );
  CIVDX1 U901 ( .A(f37[11]), .Z1(n896) );
  CNIVX1 U902 ( .A(n896), .Z(n895) );
  CIVDX1 U903 ( .A(f54[11]), .Z1(n898) );
  CNIVX1 U904 ( .A(n898), .Z(n897) );
  CIVDX1 U905 ( .A(f54[0]), .Z1(n900) );
  CNIVX1 U906 ( .A(n900), .Z(n899) );
  CIVDX1 U907 ( .A(f37[3]), .Z1(n902) );
  CNIVX1 U908 ( .A(n902), .Z(n901) );
  CIVDX1 U909 ( .A(f54[3]), .Z1(n904) );
  CNIVX1 U910 ( .A(n904), .Z(n903) );
  CIVDX1 U911 ( .A(f54[15]), .Z1(n906) );
  CNIVX1 U912 ( .A(n906), .Z(n905) );
  CIVDX1 U913 ( .A(f37[0]), .Z1(n908) );
  CNIVX1 U914 ( .A(n908), .Z(n907) );
  CIVDX1 U915 ( .A(f37[13]), .Z1(n910) );
  CNIVX1 U916 ( .A(n910), .Z(n909) );
  CIVDX1 U917 ( .A(f54[13]), .Z1(n912) );
  CNIVX1 U918 ( .A(n912), .Z(n911) );
  CIVDX1 U919 ( .A(f37[15]), .Z1(n914) );
  CNIVX1 U920 ( .A(n914), .Z(n913) );
  CIVDX1 U921 ( .A(f37[7]), .Z1(n916) );
  CNIVX1 U922 ( .A(n916), .Z(n915) );
  CIVDX1 U923 ( .A(f54[7]), .Z1(n918) );
  CNIVX1 U924 ( .A(n918), .Z(n917) );
  CIVDX1 U925 ( .A(f54[1]), .Z1(n920) );
  CNIVX1 U926 ( .A(n920), .Z(n919) );
  CIVDX1 U927 ( .A(f54[27]), .Z1(n922) );
  CNIVX1 U928 ( .A(n922), .Z(n921) );
  CIVDX1 U929 ( .A(f54[26]), .Z1(n924) );
  CNIVX1 U930 ( .A(n924), .Z(n923) );
  CIVDX1 U931 ( .A(f54[25]), .Z1(n926) );
  CNIVX1 U932 ( .A(n926), .Z(n925) );
  CIVDX1 U933 ( .A(f54[24]), .Z1(n928) );
  CNIVX1 U934 ( .A(n928), .Z(n927) );
  CIVDX1 U935 ( .A(f54[28]), .Z1(n930) );
  CNIVX1 U936 ( .A(n930), .Z(n929) );
  CIVDX1 U937 ( .A(f37[27]), .Z1(n932) );
  CNIVX1 U938 ( .A(n932), .Z(n931) );
  CIVDX1 U939 ( .A(f37[26]), .Z1(n934) );
  CNIVX1 U940 ( .A(n934), .Z(n933) );
  CIVDX1 U941 ( .A(f37[25]), .Z1(n936) );
  CNIVX1 U942 ( .A(n936), .Z(n935) );
  CIVDX1 U943 ( .A(f37[24]), .Z1(n938) );
  CNIVX1 U944 ( .A(n938), .Z(n937) );
  CIVDX1 U945 ( .A(f37[28]), .Z1(n940) );
  CNIVX1 U946 ( .A(n940), .Z(n939) );
  CNIVX1 U947 ( .A(n942), .Z(n941) );
  CNIVX1 U948 ( .A(f21[6]), .Z(n942) );
  CNIVX1 U949 ( .A(n944), .Z(n943) );
  CNIVX1 U950 ( .A(f21[10]), .Z(n944) );
  CNIVX1 U951 ( .A(n946), .Z(n945) );
  CNIVX1 U952 ( .A(f21[11]), .Z(n946) );
  CNIVX1 U953 ( .A(n948), .Z(n947) );
  CNIVX1 U954 ( .A(f21[8]), .Z(n948) );
  CNIVX1 U955 ( .A(n950), .Z(n949) );
  CNIVX1 U956 ( .A(f21[9]), .Z(n950) );
  CNIVX1 U957 ( .A(n952), .Z(n951) );
  CNIVX1 U958 ( .A(f21[15]), .Z(n952) );
  CNIVX1 U959 ( .A(n954), .Z(n953) );
  CNIVX1 U960 ( .A(f21[14]), .Z(n954) );
  CNIVX1 U961 ( .A(n956), .Z(n955) );
  CNIVX1 U962 ( .A(f02[2]), .Z(n956) );
  CNIVX1 U963 ( .A(n958), .Z(n957) );
  CNIVX1 U964 ( .A(f02[10]), .Z(n958) );
  CNIVX1 U965 ( .A(n960), .Z(n959) );
  CNIVX1 U966 ( .A(n961), .Z(n960) );
  CNIVX1 U967 ( .A(f02[5]), .Z(n961) );
  CNIVX1 U968 ( .A(n963), .Z(n962) );
  CNIVX1 U969 ( .A(f02[4]), .Z(n963) );
  CIVDX1 U970 ( .A(f61[6]), .Z1(n965) );
  CNIVX1 U971 ( .A(n965), .Z(n964) );
  CIVDX1 U972 ( .A(f61[5]), .Z1(n967) );
  CNIVX1 U973 ( .A(n967), .Z(n966) );
  CIVDX1 U974 ( .A(f61[2]), .Z1(n969) );
  CNIVX1 U975 ( .A(n969), .Z(n968) );
  CNIVX1 U976 ( .A(n971), .Z(n970) );
  CNIVX1 U977 ( .A(f02[14]), .Z(n971) );
  CNIVX1 U978 ( .A(n973), .Z(n972) );
  CNIVX1 U979 ( .A(n974), .Z(n973) );
  CNIVX1 U980 ( .A(f02[13]), .Z(n974) );
  CIVDX1 U981 ( .A(f52[18]), .Z1(n976) );
  CNIVX1 U982 ( .A(n976), .Z(n975) );
  CIVDX1 U983 ( .A(f52[6]), .Z1(n978) );
  CNIVX1 U984 ( .A(n978), .Z(n977) );
  CIVDX1 U985 ( .A(f52[2]), .Z1(n980) );
  CNIVX1 U986 ( .A(n980), .Z(n979) );
  CIVDX1 U987 ( .A(f61[22]), .Z1(n982) );
  CNIVX1 U988 ( .A(n982), .Z(n981) );
  CIVDX1 U989 ( .A(f61[18]), .Z1(n984) );
  CNIVX1 U990 ( .A(n984), .Z(n983) );
  CIVDX1 U991 ( .A(f41[18]), .Z1(n986) );
  CNIVX1 U992 ( .A(n986), .Z(n985) );
  CIVDX1 U993 ( .A(f41[6]), .Z1(n988) );
  CNIVX1 U994 ( .A(n988), .Z(n987) );
  CIVDX1 U995 ( .A(f41[2]), .Z1(n990) );
  CNIVX1 U996 ( .A(n990), .Z(n989) );
  CIVDX1 U997 ( .A(f52[22]), .Z1(n992) );
  CNIVX1 U998 ( .A(n992), .Z(n991) );
  CIVDX1 U999 ( .A(f52[20]), .Z1(n994) );
  CNIVX1 U1000 ( .A(n994), .Z(n993) );
  CIVDX1 U1001 ( .A(f31[18]), .Z1(n996) );
  CNIVX1 U1002 ( .A(n996), .Z(n995) );
  CIVDX1 U1003 ( .A(f31[6]), .Z1(n998) );
  CNIVX1 U1004 ( .A(n998), .Z(n997) );
  CIVDX1 U1005 ( .A(f31[2]), .Z1(n1000) );
  CNIVX1 U1006 ( .A(n1000), .Z(n999) );
  CIVDX1 U1007 ( .A(f41[22]), .Z1(n1002) );
  CNIVX1 U1008 ( .A(n1002), .Z(n1001) );
  CIVDX1 U1009 ( .A(f41[20]), .Z1(n1004) );
  CNIVX1 U1010 ( .A(n1004), .Z(n1003) );
  CIVDX1 U1011 ( .A(f28[18]), .Z1(n1006) );
  CNIVX1 U1012 ( .A(n1006), .Z(n1005) );
  CIVDX1 U1013 ( .A(f28[6]), .Z1(n1008) );
  CNIVX1 U1014 ( .A(n1008), .Z(n1007) );
  CIVDX1 U1015 ( .A(f28[2]), .Z1(n1010) );
  CNIVX1 U1016 ( .A(n1010), .Z(n1009) );
  CIVDX1 U1017 ( .A(f31[22]), .Z1(n1012) );
  CNIVX1 U1018 ( .A(n1012), .Z(n1011) );
  CIVDX1 U1019 ( .A(f31[20]), .Z1(n1014) );
  CNIVX1 U1020 ( .A(n1014), .Z(n1013) );
  CIVDX1 U1021 ( .A(f26[18]), .Z1(n1016) );
  CNIVX1 U1022 ( .A(n1016), .Z(n1015) );
  CIVDX1 U1023 ( .A(f26[6]), .Z1(n1018) );
  CNIVX1 U1024 ( .A(n1018), .Z(n1017) );
  CIVDX1 U1025 ( .A(f26[2]), .Z1(n1020) );
  CNIVX1 U1026 ( .A(n1020), .Z(n1019) );
  CIVDX1 U1027 ( .A(f28[22]), .Z1(n1022) );
  CNIVX1 U1028 ( .A(n1022), .Z(n1021) );
  CIVDX1 U1029 ( .A(f28[20]), .Z1(n1024) );
  CNIVX1 U1030 ( .A(n1024), .Z(n1023) );
  CIVDX1 U1031 ( .A(f28[1]), .Z1(n1026) );
  CNIVX1 U1032 ( .A(n1026), .Z(n1025) );
  CIVDX1 U1033 ( .A(f41[1]), .Z1(n1028) );
  CNIVX1 U1034 ( .A(n1028), .Z(n1027) );
  CIVDX1 U1035 ( .A(f52[1]), .Z1(n1030) );
  CNIVX1 U1036 ( .A(n1030), .Z(n1029) );
  CIVDX1 U1037 ( .A(f26[22]), .Z1(n1032) );
  CNIVX1 U1038 ( .A(n1032), .Z(n1031) );
  CIVDX1 U1039 ( .A(f26[20]), .Z1(n1034) );
  CNIVX1 U1040 ( .A(n1034), .Z(n1033) );
  CIVDX1 U1041 ( .A(f28[12]), .Z1(n1036) );
  CNIVX1 U1042 ( .A(n1036), .Z(n1035) );
  CIVDX1 U1043 ( .A(f31[12]), .Z1(n1038) );
  CNIVX1 U1044 ( .A(n1038), .Z(n1037) );
  CIVDX1 U1045 ( .A(f41[12]), .Z1(n1040) );
  CNIVX1 U1046 ( .A(n1040), .Z(n1039) );
  CIVDX1 U1047 ( .A(f52[12]), .Z1(n1042) );
  CNIVX1 U1048 ( .A(n1042), .Z(n1041) );
  CIVDX1 U1049 ( .A(f26[10]), .Z1(n1044) );
  CNIVX1 U1050 ( .A(n1044), .Z(n1043) );
  CIVDX1 U1051 ( .A(f52[7]), .Z1(n1046) );
  CNIVX1 U1052 ( .A(n1046), .Z(n1045) );
  CIVDX1 U1053 ( .A(f28[14]), .Z1(n1048) );
  CNIVX1 U1054 ( .A(n1048), .Z(n1047) );
  CIVDX1 U1055 ( .A(f31[14]), .Z1(n1050) );
  CNIVX1 U1056 ( .A(n1050), .Z(n1049) );
  CIVDX1 U1057 ( .A(f41[14]), .Z1(n1052) );
  CNIVX1 U1058 ( .A(n1052), .Z(n1051) );
  CIVDX1 U1059 ( .A(f52[14]), .Z1(n1054) );
  CNIVX1 U1060 ( .A(n1054), .Z(n1053) );
  CIVDX1 U1061 ( .A(f41[13]), .Z1(n1056) );
  CNIVX1 U1062 ( .A(n1056), .Z(n1055) );
  CIVDX1 U1063 ( .A(f52[13]), .Z1(n1058) );
  CNIVX1 U1064 ( .A(n1058), .Z(n1057) );
  CIVDX1 U1065 ( .A(f28[7]), .Z1(n1060) );
  CNIVX1 U1066 ( .A(n1060), .Z(n1059) );
  CIVDX1 U1067 ( .A(f31[7]), .Z1(n1062) );
  CNIVX1 U1068 ( .A(n1062), .Z(n1061) );
  CIVDX1 U1069 ( .A(f41[7]), .Z1(n1064) );
  CNIVX1 U1070 ( .A(n1064), .Z(n1063) );
  CIVDX1 U1071 ( .A(f31[15]), .Z1(n1066) );
  CNIVX1 U1072 ( .A(n1066), .Z(n1065) );
  CIVDX1 U1073 ( .A(f41[15]), .Z1(n1068) );
  CNIVX1 U1074 ( .A(n1068), .Z(n1067) );
  CIVDX1 U1075 ( .A(f52[15]), .Z1(n1070) );
  CNIVX1 U1076 ( .A(n1070), .Z(n1069) );
  CIVDX1 U1077 ( .A(f28[13]), .Z1(n1072) );
  CNIVX1 U1078 ( .A(n1072), .Z(n1071) );
  CIVDX1 U1079 ( .A(f31[13]), .Z1(n1074) );
  CNIVX1 U1080 ( .A(n1074), .Z(n1073) );
  CIVDX1 U1081 ( .A(f28[10]), .Z1(n1076) );
  CNIVX1 U1082 ( .A(n1076), .Z(n1075) );
  CIVDX1 U1083 ( .A(f31[10]), .Z1(n1078) );
  CNIVX1 U1084 ( .A(n1078), .Z(n1077) );
  CIVDX1 U1085 ( .A(f41[10]), .Z1(n1080) );
  CNIVX1 U1086 ( .A(n1080), .Z(n1079) );
  CIVDX1 U1087 ( .A(f52[10]), .Z1(n1082) );
  CNIVX1 U1088 ( .A(n1082), .Z(n1081) );
  CIVDX1 U1089 ( .A(f28[15]), .Z1(n1084) );
  CNIVX1 U1090 ( .A(n1084), .Z(n1083) );
  CIVDX1 U1091 ( .A(f61[9]), .Z1(n1086) );
  CNIVX1 U1092 ( .A(n1086), .Z(n1085) );
  CIVDX1 U1093 ( .A(f61[8]), .Z1(n1088) );
  CNIVX1 U1094 ( .A(n1088), .Z(n1087) );
  CIVDX1 U1095 ( .A(f61[7]), .Z1(n1090) );
  CNIVX1 U1096 ( .A(n1090), .Z(n1089) );
  CIVDX1 U1097 ( .A(f61[4]), .Z1(n1092) );
  CNIVX1 U1098 ( .A(n1092), .Z(n1091) );
  CIVDX1 U1099 ( .A(f61[0]), .Z1(n1094) );
  CNIVX1 U1100 ( .A(n1094), .Z(n1093) );
  CIVDX1 U1101 ( .A(f61[14]), .Z1(n1096) );
  CNIVX1 U1102 ( .A(n1096), .Z(n1095) );
  CIVDX1 U1103 ( .A(f61[13]), .Z1(n1098) );
  CNIVX1 U1104 ( .A(n1098), .Z(n1097) );
  CIVDX1 U1105 ( .A(f61[12]), .Z1(n1100) );
  CNIVX1 U1106 ( .A(n1100), .Z(n1099) );
  CIVDX1 U1107 ( .A(f61[11]), .Z1(n1102) );
  CNIVX1 U1108 ( .A(n1102), .Z(n1101) );
  CIVDX1 U1109 ( .A(f61[10]), .Z1(n1104) );
  CNIVX1 U1110 ( .A(n1104), .Z(n1103) );
  CIVDX1 U1111 ( .A(f61[20]), .Z1(n1106) );
  CNIVX1 U1112 ( .A(n1106), .Z(n1105) );
  CIVDX1 U1113 ( .A(f61[19]), .Z1(n1108) );
  CNIVX1 U1114 ( .A(n1108), .Z(n1107) );
  CIVDX1 U1115 ( .A(f61[17]), .Z1(n1110) );
  CNIVX1 U1116 ( .A(n1110), .Z(n1109) );
  CIVDX1 U1117 ( .A(f61[16]), .Z1(n1112) );
  CNIVX1 U1118 ( .A(n1112), .Z(n1111) );
  CIVDX1 U1119 ( .A(f61[15]), .Z1(n1114) );
  CNIVX1 U1120 ( .A(n1114), .Z(n1113) );
  CIVDX1 U1121 ( .A(f52[4]), .Z1(n1116) );
  CNIVX1 U1122 ( .A(n1116), .Z(n1115) );
  CIVDX1 U1123 ( .A(f61[25]), .Z1(n1118) );
  CNIVX1 U1124 ( .A(n1118), .Z(n1117) );
  CIVDX1 U1125 ( .A(f61[24]), .Z1(n1120) );
  CNIVX1 U1126 ( .A(n1120), .Z(n1119) );
  CIVDX1 U1127 ( .A(f61[23]), .Z1(n1122) );
  CNIVX1 U1128 ( .A(n1122), .Z(n1121) );
  CIVDX1 U1129 ( .A(f61[21]), .Z1(n1124) );
  CNIVX1 U1130 ( .A(n1124), .Z(n1123) );
  CIVDX1 U1131 ( .A(f52[19]), .Z1(n1126) );
  CNIVX1 U1132 ( .A(n1126), .Z(n1125) );
  CIVDX1 U1133 ( .A(f52[17]), .Z1(n1128) );
  CNIVX1 U1134 ( .A(n1128), .Z(n1127) );
  CIVDX1 U1135 ( .A(f52[16]), .Z1(n1130) );
  CNIVX1 U1136 ( .A(n1130), .Z(n1129) );
  CIVDX1 U1137 ( .A(f52[8]), .Z1(n1132) );
  CNIVX1 U1138 ( .A(n1132), .Z(n1131) );
  CIVDX1 U1139 ( .A(f52[5]), .Z1(n1134) );
  CNIVX1 U1140 ( .A(n1134), .Z(n1133) );
  CIVDX1 U1141 ( .A(f41[8]), .Z1(n1136) );
  CNIVX1 U1142 ( .A(n1136), .Z(n1135) );
  CIVDX1 U1143 ( .A(f41[5]), .Z1(n1138) );
  CNIVX1 U1144 ( .A(n1138), .Z(n1137) );
  CIVDX1 U1145 ( .A(f41[4]), .Z1(n1140) );
  CNIVX1 U1146 ( .A(n1140), .Z(n1139) );
  CIVDX1 U1147 ( .A(f52[23]), .Z1(n1142) );
  CNIVX1 U1148 ( .A(n1142), .Z(n1141) );
  CIVDX1 U1149 ( .A(f52[21]), .Z1(n1144) );
  CNIVX1 U1150 ( .A(n1144), .Z(n1143) );
  CIVDX1 U1151 ( .A(f41[23]), .Z1(n1146) );
  CNIVX1 U1152 ( .A(n1146), .Z(n1145) );
  CIVDX1 U1153 ( .A(f41[21]), .Z1(n1148) );
  CNIVX1 U1154 ( .A(n1148), .Z(n1147) );
  CIVDX1 U1155 ( .A(f41[19]), .Z1(n1150) );
  CNIVX1 U1156 ( .A(n1150), .Z(n1149) );
  CIVDX1 U1157 ( .A(f41[17]), .Z1(n1152) );
  CNIVX1 U1158 ( .A(n1152), .Z(n1151) );
  CIVDX1 U1159 ( .A(f41[16]), .Z1(n1154) );
  CNIVX1 U1160 ( .A(n1154), .Z(n1153) );
  CIVDX1 U1161 ( .A(f31[17]), .Z1(n1156) );
  CNIVX1 U1162 ( .A(n1156), .Z(n1155) );
  CIVDX1 U1163 ( .A(f31[16]), .Z1(n1158) );
  CNIVX1 U1164 ( .A(n1158), .Z(n1157) );
  CIVDX1 U1165 ( .A(f31[8]), .Z1(n1160) );
  CNIVX1 U1166 ( .A(n1160), .Z(n1159) );
  CIVDX1 U1167 ( .A(f31[5]), .Z1(n1162) );
  CNIVX1 U1168 ( .A(n1162), .Z(n1161) );
  CIVDX1 U1169 ( .A(f31[4]), .Z1(n1164) );
  CNIVX1 U1170 ( .A(n1164), .Z(n1163) );
  CIVDX1 U1171 ( .A(f28[5]), .Z1(n1166) );
  CNIVX1 U1172 ( .A(n1166), .Z(n1165) );
  CIVDX1 U1173 ( .A(f28[4]), .Z1(n1168) );
  CNIVX1 U1174 ( .A(n1168), .Z(n1167) );
  CIVDX1 U1175 ( .A(f31[23]), .Z1(n1170) );
  CNIVX1 U1176 ( .A(n1170), .Z(n1169) );
  CIVDX1 U1177 ( .A(f31[21]), .Z1(n1172) );
  CNIVX1 U1178 ( .A(n1172), .Z(n1171) );
  CIVDX1 U1179 ( .A(f31[19]), .Z1(n1174) );
  CNIVX1 U1180 ( .A(n1174), .Z(n1173) );
  CIVDX1 U1181 ( .A(f28[21]), .Z1(n1176) );
  CNIVX1 U1182 ( .A(n1176), .Z(n1175) );
  CIVDX1 U1183 ( .A(f28[19]), .Z1(n1178) );
  CNIVX1 U1184 ( .A(n1178), .Z(n1177) );
  CIVDX1 U1185 ( .A(f28[17]), .Z1(n1180) );
  CNIVX1 U1186 ( .A(n1180), .Z(n1179) );
  CIVDX1 U1187 ( .A(f28[16]), .Z1(n1182) );
  CNIVX1 U1188 ( .A(n1182), .Z(n1181) );
  CIVDX1 U1189 ( .A(f28[8]), .Z1(n1184) );
  CNIVX1 U1190 ( .A(n1184), .Z(n1183) );
  CIVDX1 U1191 ( .A(f26[8]), .Z1(n1186) );
  CNIVX1 U1192 ( .A(n1186), .Z(n1185) );
  CIVDX1 U1193 ( .A(f26[7]), .Z1(n1188) );
  CNIVX1 U1194 ( .A(n1188), .Z(n1187) );
  CIVDX1 U1195 ( .A(f26[5]), .Z1(n1190) );
  CNIVX1 U1196 ( .A(n1190), .Z(n1189) );
  CIVDX1 U1197 ( .A(f26[4]), .Z1(n1192) );
  CNIVX1 U1198 ( .A(n1192), .Z(n1191) );
  CIVDX1 U1199 ( .A(f28[23]), .Z1(n1194) );
  CNIVX1 U1200 ( .A(n1194), .Z(n1193) );
  CIVDX1 U1201 ( .A(f26[16]), .Z1(n1196) );
  CNIVX1 U1202 ( .A(n1196), .Z(n1195) );
  CIVDX1 U1203 ( .A(f26[15]), .Z1(n1198) );
  CNIVX1 U1204 ( .A(n1198), .Z(n1197) );
  CIVDX1 U1205 ( .A(f26[14]), .Z1(n1200) );
  CNIVX1 U1206 ( .A(n1200), .Z(n1199) );
  CIVDX1 U1207 ( .A(f26[13]), .Z1(n1202) );
  CNIVX1 U1208 ( .A(n1202), .Z(n1201) );
  CIVDX1 U1209 ( .A(f26[12]), .Z1(n1204) );
  CNIVX1 U1210 ( .A(n1204), .Z(n1203) );
  CIVDX1 U1211 ( .A(f61[1]), .Z1(n1206) );
  CNIVX1 U1212 ( .A(n1206), .Z(n1205) );
  CIVDX1 U1213 ( .A(f26[23]), .Z1(n1208) );
  CNIVX1 U1214 ( .A(n1208), .Z(n1207) );
  CIVDX1 U1215 ( .A(f26[21]), .Z1(n1210) );
  CNIVX1 U1216 ( .A(n1210), .Z(n1209) );
  CIVDX1 U1217 ( .A(f26[19]), .Z1(n1212) );
  CNIVX1 U1218 ( .A(n1212), .Z(n1211) );
  CIVDX1 U1219 ( .A(f26[17]), .Z1(n1214) );
  CNIVX1 U1220 ( .A(n1214), .Z(n1213) );
  CIVDX1 U1221 ( .A(f31[3]), .Z1(n1216) );
  CNIVX1 U1222 ( .A(n1216), .Z(n1215) );
  CIVDX1 U1223 ( .A(f41[3]), .Z1(n1218) );
  CNIVX1 U1224 ( .A(n1218), .Z(n1217) );
  CIVDX1 U1225 ( .A(f52[3]), .Z1(n1220) );
  CNIVX1 U1226 ( .A(n1220), .Z(n1219) );
  CIVDX1 U1227 ( .A(f26[1]), .Z1(n1222) );
  CNIVX1 U1228 ( .A(n1222), .Z(n1221) );
  CIVDX1 U1229 ( .A(f61[3]), .Z1(n1224) );
  CNIVX1 U1230 ( .A(n1224), .Z(n1223) );
  CIVDX1 U1231 ( .A(f28[9]), .Z1(n1226) );
  CNIVX1 U1232 ( .A(n1226), .Z(n1225) );
  CIVDX1 U1233 ( .A(f31[9]), .Z1(n1228) );
  CNIVX1 U1234 ( .A(n1228), .Z(n1227) );
  CIVDX1 U1235 ( .A(f41[9]), .Z1(n1230) );
  CNIVX1 U1236 ( .A(n1230), .Z(n1229) );
  CIVDX1 U1237 ( .A(f52[9]), .Z1(n1232) );
  CNIVX1 U1238 ( .A(n1232), .Z(n1231) );
  CIVDX1 U1239 ( .A(f28[3]), .Z1(n1234) );
  CNIVX1 U1240 ( .A(n1234), .Z(n1233) );
  CIVDX1 U1241 ( .A(f26[3]), .Z1(n1236) );
  CNIVX1 U1242 ( .A(n1236), .Z(n1235) );
  CIVDX1 U1243 ( .A(f28[11]), .Z1(n1238) );
  CNIVX1 U1244 ( .A(n1238), .Z(n1237) );
  CIVDX1 U1245 ( .A(f31[11]), .Z1(n1240) );
  CNIVX1 U1246 ( .A(n1240), .Z(n1239) );
  CIVDX1 U1247 ( .A(f41[11]), .Z1(n1242) );
  CNIVX1 U1248 ( .A(n1242), .Z(n1241) );
  CIVDX1 U1249 ( .A(f52[11]), .Z1(n1244) );
  CNIVX1 U1250 ( .A(n1244), .Z(n1243) );
  CIVDX1 U1251 ( .A(f26[0]), .Z1(n1246) );
  CNIVX1 U1252 ( .A(n1246), .Z(n1245) );
  CIVDX1 U1253 ( .A(f28[0]), .Z1(n1248) );
  CNIVX1 U1254 ( .A(n1248), .Z(n1247) );
  CIVDX1 U1255 ( .A(f31[0]), .Z1(n1250) );
  CNIVX1 U1256 ( .A(n1250), .Z(n1249) );
  CIVDX1 U1257 ( .A(f41[0]), .Z1(n1252) );
  CNIVX1 U1258 ( .A(n1252), .Z(n1251) );
  CIVDX1 U1259 ( .A(f52[0]), .Z1(n1254) );
  CNIVX1 U1260 ( .A(n1254), .Z(n1253) );
  CIVDX1 U1261 ( .A(f61[28]), .Z1(n1256) );
  CNIVX1 U1262 ( .A(n1256), .Z(n1255) );
  CIVDX1 U1263 ( .A(f61[27]), .Z1(n1258) );
  CNIVX1 U1264 ( .A(n1258), .Z(n1257) );
  CIVDX1 U1265 ( .A(f61[26]), .Z1(n1260) );
  CNIVX1 U1266 ( .A(n1260), .Z(n1259) );
  CIVDX1 U1267 ( .A(f26[9]), .Z1(n1262) );
  CNIVX1 U1268 ( .A(n1262), .Z(n1261) );
  CIVDX1 U1269 ( .A(f26[11]), .Z1(n1264) );
  CNIVX1 U1270 ( .A(n1264), .Z(n1263) );
  CIVDX1 U1271 ( .A(f52[28]), .Z1(n1266) );
  CNIVX1 U1272 ( .A(n1266), .Z(n1265) );
  CIVDX1 U1273 ( .A(f52[27]), .Z1(n1268) );
  CNIVX1 U1274 ( .A(n1268), .Z(n1267) );
  CIVDX1 U1275 ( .A(f52[26]), .Z1(n1270) );
  CNIVX1 U1276 ( .A(n1270), .Z(n1269) );
  CIVDX1 U1277 ( .A(f52[25]), .Z1(n1272) );
  CNIVX1 U1278 ( .A(n1272), .Z(n1271) );
  CIVDX1 U1279 ( .A(f52[24]), .Z1(n1274) );
  CNIVX1 U1280 ( .A(n1274), .Z(n1273) );
  CIVDX1 U1281 ( .A(f41[28]), .Z1(n1276) );
  CNIVX1 U1282 ( .A(n1276), .Z(n1275) );
  CIVDX1 U1283 ( .A(f41[27]), .Z1(n1278) );
  CNIVX1 U1284 ( .A(n1278), .Z(n1277) );
  CIVDX1 U1285 ( .A(f41[26]), .Z1(n1280) );
  CNIVX1 U1286 ( .A(n1280), .Z(n1279) );
  CIVDX1 U1287 ( .A(f41[25]), .Z1(n1282) );
  CNIVX1 U1288 ( .A(n1282), .Z(n1281) );
  CIVDX1 U1289 ( .A(f41[24]), .Z1(n1284) );
  CNIVX1 U1290 ( .A(n1284), .Z(n1283) );
  CIVDX1 U1291 ( .A(f31[28]), .Z1(n1286) );
  CNIVX1 U1292 ( .A(n1286), .Z(n1285) );
  CIVDX1 U1293 ( .A(f31[27]), .Z1(n1288) );
  CNIVX1 U1294 ( .A(n1288), .Z(n1287) );
  CIVDX1 U1295 ( .A(f31[26]), .Z1(n1290) );
  CNIVX1 U1296 ( .A(n1290), .Z(n1289) );
  CIVDX1 U1297 ( .A(f31[25]), .Z1(n1292) );
  CNIVX1 U1298 ( .A(n1292), .Z(n1291) );
  CIVDX1 U1299 ( .A(f31[24]), .Z1(n1294) );
  CNIVX1 U1300 ( .A(n1294), .Z(n1293) );
  CIVDX1 U1301 ( .A(f28[28]), .Z1(n1296) );
  CNIVX1 U1302 ( .A(n1296), .Z(n1295) );
  CIVDX1 U1303 ( .A(f28[27]), .Z1(n1298) );
  CNIVX1 U1304 ( .A(n1298), .Z(n1297) );
  CIVDX1 U1305 ( .A(f28[26]), .Z1(n1300) );
  CNIVX1 U1306 ( .A(n1300), .Z(n1299) );
  CIVDX1 U1307 ( .A(f28[25]), .Z1(n1302) );
  CNIVX1 U1308 ( .A(n1302), .Z(n1301) );
  CIVDX1 U1309 ( .A(f28[24]), .Z1(n1304) );
  CNIVX1 U1310 ( .A(n1304), .Z(n1303) );
  CIVDX1 U1311 ( .A(f26[28]), .Z1(n1306) );
  CNIVX1 U1312 ( .A(n1306), .Z(n1305) );
  CIVDX1 U1313 ( .A(f26[27]), .Z1(n1308) );
  CNIVX1 U1314 ( .A(n1308), .Z(n1307) );
  CIVDX1 U1315 ( .A(f26[26]), .Z1(n1310) );
  CNIVX1 U1316 ( .A(n1310), .Z(n1309) );
  CIVDX1 U1317 ( .A(f26[25]), .Z1(n1312) );
  CNIVX1 U1318 ( .A(n1312), .Z(n1311) );
  CIVDX1 U1319 ( .A(f26[24]), .Z1(n1314) );
  CNIVX1 U1320 ( .A(n1314), .Z(n1313) );
  CNIVX1 U1321 ( .A(f02[30]), .Z(n1315) );
  CNIVX1 U1322 ( .A(n1317), .Z(n1316) );
  CNIVX1 U1323 ( .A(captA[25]), .Z(n1317) );
  CNIVX1 U1324 ( .A(f01[29]), .Z(n1318) );
  CNIVX1 U1325 ( .A(f01[28]), .Z(n1319) );
  CIVDX1 U1326 ( .A(f31[1]), .Z1(n1321) );
  CNIVX1 U1327 ( .A(n1321), .Z(n1320) );
  CNIVX1 U1328 ( .A(f01[30]), .Z(n1322) );
  CNIVX1 U1329 ( .A(n1324), .Z(n1323) );
  CNIVX1 U1330 ( .A(f11[31]), .Z(n1324) );
  CNIVX1 U1331 ( .A(n1326), .Z(n1325) );
  CNIVX1 U1332 ( .A(f11[30]), .Z(n1326) );
  CMX2X1 U1333 ( .A0(f27[25]), .A1(f38[25]), .S(rst), .Z(n79) );
  CNIVX2 U1334 ( .A(f21[29]), .Z(n1327) );
  CIVDX1 U1335 ( .A(f37[29]), .Z1(n1329) );
  CNIVX1 U1336 ( .A(n1329), .Z(n1328) );
  CIVDX1 U1337 ( .A(f54[29]), .Z1(n1331) );
  CNIVX1 U1338 ( .A(n1331), .Z(n1330) );
  CIVDX1 U1339 ( .A(f37[31]), .Z1(n1333) );
  CNIVX1 U1340 ( .A(n1333), .Z(n1332) );
  CIVDX1 U1341 ( .A(f54[31]), .Z1(n1335) );
  CNIVX1 U1342 ( .A(n1335), .Z(n1334) );
  CIVDX1 U1343 ( .A(f41[29]), .Z1(n1337) );
  CNIVX1 U1344 ( .A(n1337), .Z(n1336) );
  CIVDX1 U1345 ( .A(f52[29]), .Z1(n1339) );
  CNIVX1 U1346 ( .A(n1339), .Z(n1338) );
  CIVDX1 U1347 ( .A(f61[30]), .Z1(n1341) );
  CNIVX1 U1348 ( .A(n1341), .Z(n1340) );
  CIVDX1 U1349 ( .A(f61[29]), .Z1(n1343) );
  CNIVX1 U1350 ( .A(n1343), .Z(n1342) );
  CIVDX1 U1351 ( .A(f52[31]), .Z1(n1345) );
  CNIVX1 U1352 ( .A(n1345), .Z(n1344) );
  CIVDX1 U1353 ( .A(f61[31]), .Z1(n1347) );
  CNIVX1 U1354 ( .A(n1347), .Z(n1346) );
  CIVDX1 U1355 ( .A(f26[29]), .Z1(n1349) );
  CNIVX1 U1356 ( .A(n1349), .Z(n1348) );
  CIVDX1 U1357 ( .A(f28[29]), .Z1(n1351) );
  CNIVX1 U1358 ( .A(n1351), .Z(n1350) );
  CIVDX1 U1359 ( .A(f31[29]), .Z1(n1353) );
  CNIVX1 U1360 ( .A(n1353), .Z(n1352) );
  CNIVX1 U1361 ( .A(n1355), .Z(n1354) );
  CNIVX1 U1362 ( .A(f21[30]), .Z(n1355) );
  CIVDX1 U1363 ( .A(f26[31]), .Z1(n1357) );
  CNIVX1 U1364 ( .A(n1357), .Z(n1356) );
  CIVDX1 U1365 ( .A(f28[31]), .Z1(n1359) );
  CNIVX1 U1366 ( .A(n1359), .Z(n1358) );
  CIVDX1 U1367 ( .A(f31[31]), .Z1(n1361) );
  CNIVX1 U1368 ( .A(n1361), .Z(n1360) );
  CIVDX1 U1369 ( .A(f41[31]), .Z1(n1363) );
  CNIVX1 U1370 ( .A(n1363), .Z(n1362) );
  CIVDX1 U1371 ( .A(f37[30]), .Z1(n1365) );
  CNIVX1 U1372 ( .A(n1365), .Z(n1364) );
  CIVDX1 U1373 ( .A(f54[30]), .Z1(n1367) );
  CNIVX1 U1374 ( .A(n1367), .Z(n1366) );
  CIVDX1 U1375 ( .A(f26[30]), .Z1(n1369) );
  CNIVX1 U1376 ( .A(n1369), .Z(n1368) );
  CIVDX1 U1377 ( .A(f28[30]), .Z1(n1371) );
  CNIVX1 U1378 ( .A(n1371), .Z(n1370) );
  CIVDX1 U1379 ( .A(n1418), .Z1(n1373) );
  CNIVX1 U1380 ( .A(n1373), .Z(n1372) );
  CIVDX1 U1381 ( .A(f41[30]), .Z1(n1375) );
  CNIVX1 U1382 ( .A(n1375), .Z(n1374) );
  CIVDX1 U1383 ( .A(f52[30]), .Z1(n1377) );
  CNIVX1 U1384 ( .A(n1377), .Z(n1376) );
  CNIVX1 U1385 ( .A(n1516), .Z(n1381) );
  CNIVX1 U1386 ( .A(n1383), .Z(n1382) );
  CNIVX1 U1387 ( .A(f21[31]), .Z(n1383) );
  CNIVX1 U1388 ( .A(res_d[30]), .Z(n1384) );
  CNIVX1 U1389 ( .A(res_d[31]), .Z(n1385) );
  CNIVX1 U1390 ( .A(res_d[25]), .Z(n1386) );
  CNIVX1 U1391 ( .A(res_d[26]), .Z(n1387) );
  CNIVX1 U1392 ( .A(res_d[27]), .Z(n1388) );
  CNIVX1 U1393 ( .A(res_d[28]), .Z(n1389) );
  CNIVX1 U1394 ( .A(res_d[29]), .Z(n1390) );
  CNIVX1 U1395 ( .A(res_d[20]), .Z(n1391) );
  CNIVX1 U1396 ( .A(res_d[21]), .Z(n1392) );
  CNIVX1 U1397 ( .A(res_d[22]), .Z(n1393) );
  CNIVX1 U1398 ( .A(res_d[23]), .Z(n1394) );
  CNIVX1 U1399 ( .A(res_d[24]), .Z(n1395) );
  CNIVX1 U1400 ( .A(res_d[15]), .Z(n1396) );
  CNIVX1 U1401 ( .A(res_d[16]), .Z(n1397) );
  CNIVX1 U1402 ( .A(res_d[17]), .Z(n1398) );
  CNIVX1 U1403 ( .A(res_d[18]), .Z(n1399) );
  CNIVX1 U1404 ( .A(res_d[19]), .Z(n1400) );
  CNIVX1 U1405 ( .A(res_d[10]), .Z(n1401) );
  CNIVX1 U1406 ( .A(res_d[11]), .Z(n1402) );
  CNIVX1 U1407 ( .A(res_d[12]), .Z(n1403) );
  CNIVX1 U1408 ( .A(res_d[13]), .Z(n1404) );
  CNIVX1 U1409 ( .A(res_d[14]), .Z(n1405) );
  CNIVX1 U1410 ( .A(res_d[5]), .Z(n1406) );
  CNIVX1 U1411 ( .A(res_d[6]), .Z(n1407) );
  CNIVX1 U1412 ( .A(res_d[7]), .Z(n1408) );
  CNIVX1 U1413 ( .A(res_d[8]), .Z(n1409) );
  CNIVX1 U1414 ( .A(res_d[9]), .Z(n1410) );
  CNIVX1 U1415 ( .A(res_d[0]), .Z(n1411) );
  CNIVX1 U1416 ( .A(res_d[1]), .Z(n1412) );
  CNIVX1 U1417 ( .A(res_d[2]), .Z(n1413) );
  CNIVX1 U1418 ( .A(res_d[3]), .Z(n1414) );
  CNIVX1 U1419 ( .A(res_d[4]), .Z(n1415) );
  CIVX2 U1420 ( .A(w5[17]), .Z(n1416) );
  CIVX4 U1421 ( .A(n1416), .Z(n1417) );
  CMX2XL U1422 ( .A0(n332), .A1(C[17]), .S(n18), .Z(n103) );
  CMX2XL U1423 ( .A0(n272), .A1(B[2]), .S(n20), .Z(n120) );
  CMX2XL U1424 ( .A0(n443), .A1(A[2]), .S(n16), .Z(n152) );
  CMX2XL U1425 ( .A0(n481), .A1(C[2]), .S(n18), .Z(n88) );
  CNIVX2 U1426 ( .A(w5[24]), .Z(n1421) );
  CNR2XL U1427 ( .A(stopB), .B(pushB), .Z(n14) );
  CNR2XL U1428 ( .A(pushA), .B(stopA), .Z(n13) );
  CNR2XL U1429 ( .A(pushC), .B(stopC), .Z(n15) );
  CMX2XL U1430 ( .A0(captC[28]), .A1(C[28]), .S(n18), .Z(n114) );
  CMX2XL U1431 ( .A0(captC[30]), .A1(C[30]), .S(n18), .Z(n116) );
  CMX2XL U1432 ( .A0(captB[28]), .A1(B[28]), .S(n20), .Z(n146) );
  CMX2XL U1433 ( .A0(captB[30]), .A1(B[30]), .S(n20), .Z(n148) );
  CMX2XL U1434 ( .A0(captA[28]), .A1(A[28]), .S(n16), .Z(n178) );
  CMX2XL U1435 ( .A0(captA[30]), .A1(A[30]), .S(n16), .Z(n180) );
  CAOR2XL U1436 ( .A(C[31]), .B(n18), .C(n1380), .D(n1526), .Z(n117) );
  CAOR2XL U1437 ( .A(B[31]), .B(n20), .C(n1379), .D(n1525), .Z(n149) );
  CAOR2XL U1438 ( .A(A[31]), .B(n16), .C(n1378), .D(n1524), .Z(n181) );
  CNR3XL U1439 ( .A(n15), .B(n13), .C(n14), .Z(N7) );
  CIVX2 U1440 ( .A(n1526), .Z(n18) );
  CIVX2 U1441 ( .A(n1525), .Z(n20) );
  CIVX2 U1442 ( .A(n1524), .Z(n16) );
  CNR2X1 U1443 ( .A(N7), .B(n14), .Z(seen_d[1]) );
  CNR2X1 U1444 ( .A(N7), .B(n13), .Z(seen_d[2]) );
  CNR2X1 U1445 ( .A(N7), .B(n15), .Z(seen_d[0]) );
  CNIVX1 U1446 ( .A(n1513), .Z(n1424) );
  CNIVX1 U1447 ( .A(n1513), .Z(n1501) );
  CNIVX1 U1448 ( .A(n1513), .Z(n1436) );
  CNIVX1 U1449 ( .A(n1513), .Z(n1493) );
  CNIVX1 U1450 ( .A(n1513), .Z(n1476) );
  CNIVX1 U1451 ( .A(n1513), .Z(n1473) );
  CNIVX1 U1452 ( .A(n1513), .Z(n1498) );
  CNIVX1 U1453 ( .A(n1513), .Z(n1506) );
  CNIVX1 U1454 ( .A(n1513), .Z(n1489) );
  CNIVX1 U1455 ( .A(n1513), .Z(n1487) );
  CNIVX1 U1456 ( .A(n1513), .Z(n1484) );
  CNIVX1 U1457 ( .A(n1513), .Z(n1441) );
  CNIVX1 U1458 ( .A(n1513), .Z(n1438) );
  CNIVX1 U1459 ( .A(n1513), .Z(n1495) );
  CNIVX1 U1460 ( .A(n1513), .Z(n1509) );
  CNIVX1 U1461 ( .A(n1513), .Z(n1503) );
  CNIVX1 U1462 ( .A(n1513), .Z(n1478) );
  CNIVX1 U1463 ( .A(n1513), .Z(n1470) );
  CNIVX1 U1464 ( .A(n1513), .Z(n1481) );
  CNIVX1 U1465 ( .A(n1513), .Z(n1456) );
  CNIVX1 U1466 ( .A(n1513), .Z(n1455) );
  CNIVX1 U1467 ( .A(n1513), .Z(n1454) );
  CNIVX1 U1468 ( .A(n1513), .Z(n1453) );
  CNIVX1 U1469 ( .A(n1513), .Z(n1452) );
  CNIVX1 U1470 ( .A(n1513), .Z(n1451) );
  CNIVX1 U1471 ( .A(n1513), .Z(n1450) );
  CNIVX1 U1472 ( .A(n1513), .Z(n1449) );
  CNIVX1 U1473 ( .A(n1513), .Z(n1448) );
  CNIVX1 U1474 ( .A(n1513), .Z(n1447) );
  CNIVX1 U1475 ( .A(n1513), .Z(n1446) );
  CNIVX1 U1476 ( .A(n1513), .Z(n1467) );
  CNIVX1 U1477 ( .A(n1513), .Z(n1466) );
  CNIVX1 U1478 ( .A(n1513), .Z(n1465) );
  CNIVX1 U1479 ( .A(n1513), .Z(n1440) );
  CNIVX1 U1480 ( .A(n1513), .Z(n1439) );
  CNIVX1 U1481 ( .A(n1513), .Z(n1437) );
  CNIVX1 U1482 ( .A(n1513), .Z(n1500) );
  CNIVX1 U1483 ( .A(n1513), .Z(n1499) );
  CNIVX1 U1484 ( .A(n1513), .Z(n1497) );
  CNIVX1 U1485 ( .A(n1513), .Z(n1496) );
  CNIVX1 U1486 ( .A(n1513), .Z(n1494) );
  CNIVX1 U1487 ( .A(n1513), .Z(n1492) );
  CNIVX1 U1488 ( .A(n1513), .Z(n1491) );
  CNIVX1 U1489 ( .A(n1513), .Z(n1508) );
  CNIVX1 U1490 ( .A(n1513), .Z(n1507) );
  CNIVX1 U1491 ( .A(n1513), .Z(n1505) );
  CNIVX1 U1492 ( .A(n1513), .Z(n1504) );
  CNIVX1 U1493 ( .A(n1513), .Z(n1502) );
  CNIVX1 U1494 ( .A(n1513), .Z(n1479) );
  CNIVX1 U1495 ( .A(n1513), .Z(n1477) );
  CNIVX1 U1496 ( .A(n1513), .Z(n1475) );
  CNIVX1 U1497 ( .A(n1513), .Z(n1474) );
  CNIVX1 U1498 ( .A(n1513), .Z(n1472) );
  CNIVX1 U1499 ( .A(n1513), .Z(n1471) );
  CNIVX1 U1500 ( .A(n1513), .Z(n1469) );
  CNIVX1 U1501 ( .A(n1513), .Z(n1490) );
  CNIVX1 U1502 ( .A(n1513), .Z(n1488) );
  CNIVX1 U1503 ( .A(n1513), .Z(n1486) );
  CNIVX1 U1504 ( .A(n1513), .Z(n1485) );
  CNIVX1 U1505 ( .A(n1513), .Z(n1483) );
  CNIVX1 U1506 ( .A(n1513), .Z(n1482) );
  CNIVX1 U1507 ( .A(n1513), .Z(n1480) );
  CNIVX1 U1508 ( .A(n1513), .Z(n1462) );
  CNIVX1 U1509 ( .A(n1513), .Z(n1461) );
  CNIVX1 U1510 ( .A(n1513), .Z(n1460) );
  CNIVX1 U1511 ( .A(n1513), .Z(n1459) );
  CNIVX1 U1512 ( .A(n1513), .Z(n1458) );
  CNIVX1 U1513 ( .A(n1513), .Z(n1457) );
  CNIVX1 U1514 ( .A(n1513), .Z(n1435) );
  CNIVX1 U1515 ( .A(n1513), .Z(n1434) );
  CNIVX1 U1516 ( .A(n1513), .Z(n1433) );
  CNIVX1 U1517 ( .A(n1513), .Z(n1432) );
  CNIVX1 U1518 ( .A(n1513), .Z(n1431) );
  CNIVX1 U1519 ( .A(n1513), .Z(n1430) );
  CNIVX1 U1520 ( .A(n1513), .Z(n1429) );
  CNIVX1 U1521 ( .A(n1513), .Z(n1428) );
  CNIVX1 U1522 ( .A(n1513), .Z(n1427) );
  CNIVX1 U1523 ( .A(n1513), .Z(n1426) );
  CNIVX1 U1524 ( .A(n1513), .Z(n1425) );
  CNIVX1 U1525 ( .A(n1513), .Z(n1445) );
  CNIVX1 U1526 ( .A(n1513), .Z(n1444) );
  CNIVX1 U1527 ( .A(n1513), .Z(n1443) );
  CNIVX1 U1528 ( .A(n1513), .Z(n1442) );
  CNIVX1 U1529 ( .A(n1513), .Z(n1463) );
  CNIVX1 U1530 ( .A(n1513), .Z(n1464) );
  CNIVX1 U1531 ( .A(n1513), .Z(n1468) );
  CNIVX1 U1532 ( .A(n1513), .Z(n1510) );
  CNIVX1 U1533 ( .A(n1513), .Z(n1511) );
  CNIVX1 U1534 ( .A(n1513), .Z(n1512) );
  CNIVXL U1535 ( .A(f12[3]), .Z(n1518) );
  CNIVX1 U1536 ( .A(w5[8]), .Z(n1516) );
  CIVX2 U1541 ( .A(rst), .Z(n1513) );
  CIVXL U1542 ( .A(f12[9]), .Z(n1514) );
  CIVXL U1543 ( .A(f12[2]), .Z(n1519) );
  CIVX2 U1544 ( .A(n1519), .Z(n1520) );
  CIVX2 U1545 ( .A(stopA), .Z(n1521) );
  CND2X1 U1546 ( .A(pushA), .B(n1521), .Z(n1524) );
  CMX2X1 U1547 ( .A0(n504), .A1(A[0]), .S(n16), .Z(n150) );
  CMX2X1 U1548 ( .A0(n712), .A1(A[1]), .S(n16), .Z(n151) );
  CMX2X1 U1549 ( .A0(n708), .A1(A[3]), .S(n16), .Z(n153) );
  CMX2X1 U1550 ( .A0(n523), .A1(A[4]), .S(n16), .Z(n154) );
  CMX2X1 U1551 ( .A0(n500), .A1(A[5]), .S(n16), .Z(n155) );
  CMX2X1 U1552 ( .A0(n458), .A1(A[6]), .S(n16), .Z(n156) );
  CMX2X1 U1553 ( .A0(n486), .A1(A[7]), .S(n16), .Z(n157) );
  CMX2X1 U1554 ( .A0(n455), .A1(A[8]), .S(n16), .Z(n158) );
  CMX2X1 U1555 ( .A0(n453), .A1(A[9]), .S(n16), .Z(n159) );
  CMX2X1 U1556 ( .A0(n533), .A1(A[10]), .S(n16), .Z(n160) );
  CMX2X1 U1557 ( .A0(n518), .A1(A[11]), .S(n16), .Z(n161) );
  CMX2X1 U1558 ( .A0(n517), .A1(A[12]), .S(n16), .Z(n162) );
  CMX2X1 U1559 ( .A0(n520), .A1(A[13]), .S(n16), .Z(n163) );
  CMX2X1 U1560 ( .A0(n325), .A1(A[14]), .S(n16), .Z(n164) );
  CMX2X1 U1561 ( .A0(n519), .A1(A[15]), .S(n16), .Z(n165) );
  CMX2X1 U1562 ( .A0(n530), .A1(A[16]), .S(n16), .Z(n166) );
  CMX2X1 U1563 ( .A0(captA[17]), .A1(A[17]), .S(n16), .Z(n167) );
  CMX2X1 U1564 ( .A0(n735), .A1(A[18]), .S(n16), .Z(n168) );
  CMX2X1 U1565 ( .A0(n498), .A1(A[19]), .S(n16), .Z(n169) );
  CMX2X1 U1566 ( .A0(n248), .A1(A[20]), .S(n16), .Z(n170) );
  CMX2X1 U1567 ( .A0(captA[21]), .A1(A[21]), .S(n16), .Z(n171) );
  CMX2X1 U1568 ( .A0(captA[22]), .A1(A[22]), .S(n16), .Z(n172) );
  CMX2X1 U1569 ( .A0(captA[23]), .A1(A[23]), .S(n16), .Z(n173) );
  CMX2X1 U1570 ( .A0(captA[24]), .A1(A[24]), .S(n16), .Z(n174) );
  CMX2X1 U1571 ( .A0(captA[25]), .A1(A[25]), .S(n16), .Z(n175) );
  CMX2X1 U1572 ( .A0(captA[26]), .A1(A[26]), .S(n16), .Z(n176) );
  CMX2X1 U1573 ( .A0(captA[27]), .A1(A[27]), .S(n16), .Z(n177) );
  CMX2X1 U1574 ( .A0(captA[29]), .A1(A[29]), .S(n16), .Z(n179) );
  CIVX2 U1575 ( .A(stopB), .Z(n1522) );
  CND2X1 U1576 ( .A(pushB), .B(n1522), .Z(n1525) );
  CMX2X1 U1577 ( .A0(n681), .A1(B[0]), .S(n20), .Z(n118) );
  CMX2X1 U1578 ( .A0(n711), .A1(B[1]), .S(n20), .Z(n119) );
  CMX2X1 U1579 ( .A0(n515), .A1(B[3]), .S(n20), .Z(n121) );
  CMX2X1 U1580 ( .A0(n228), .A1(B[4]), .S(n20), .Z(n122) );
  CMX2X1 U1581 ( .A0(n683), .A1(B[5]), .S(n20), .Z(n123) );
  CMX2X1 U1582 ( .A0(n448), .A1(B[6]), .S(n20), .Z(n124) );
  CMX2X1 U1583 ( .A0(n488), .A1(B[7]), .S(n20), .Z(n125) );
  CMX2X1 U1584 ( .A0(n492), .A1(B[8]), .S(n20), .Z(n126) );
  CMX2X1 U1585 ( .A0(n363), .A1(B[9]), .S(n20), .Z(n127) );
  CMX2X1 U1586 ( .A0(captB[10]), .A1(B[10]), .S(n20), .Z(n128) );
  CMX2X1 U1587 ( .A0(n516), .A1(B[11]), .S(n20), .Z(n129) );
  CMX2X1 U1588 ( .A0(n687), .A1(B[12]), .S(n20), .Z(n130) );
  CMX2X1 U1589 ( .A0(n521), .A1(B[13]), .S(n20), .Z(n131) );
  CMX2X1 U1590 ( .A0(n514), .A1(B[14]), .S(n20), .Z(n132) );
  CMX2X1 U1591 ( .A0(n690), .A1(B[15]), .S(n20), .Z(n133) );
  CMX2X1 U1592 ( .A0(n693), .A1(B[16]), .S(n20), .Z(n134) );
  CMX2X1 U1593 ( .A0(n202), .A1(B[17]), .S(n20), .Z(n135) );
  CMX2X1 U1594 ( .A0(n696), .A1(B[18]), .S(n20), .Z(n136) );
  CMX2X1 U1595 ( .A0(n699), .A1(B[19]), .S(n20), .Z(n137) );
  CMX2X1 U1596 ( .A0(n702), .A1(B[20]), .S(n20), .Z(n138) );
  CMX2X1 U1597 ( .A0(captB[21]), .A1(B[21]), .S(n20), .Z(n139) );
  CMX2X1 U1598 ( .A0(captB[22]), .A1(B[22]), .S(n20), .Z(n140) );
  CMX2X1 U1599 ( .A0(captB[23]), .A1(B[23]), .S(n20), .Z(n141) );
  CMX2X1 U1600 ( .A0(captB[24]), .A1(B[24]), .S(n20), .Z(n142) );
  CMX2X1 U1601 ( .A0(captB[25]), .A1(B[25]), .S(n20), .Z(n143) );
  CMX2X1 U1602 ( .A0(captB[26]), .A1(B[26]), .S(n20), .Z(n144) );
  CMX2X1 U1603 ( .A0(captB[27]), .A1(B[27]), .S(n20), .Z(n145) );
  CMX2X1 U1604 ( .A0(captB[29]), .A1(B[29]), .S(n20), .Z(n147) );
  CIVX2 U1605 ( .A(stopC), .Z(n1523) );
  CND2X1 U1606 ( .A(pushC), .B(n1523), .Z(n1526) );
  CMX2X1 U1607 ( .A0(n527), .A1(C[0]), .S(n18), .Z(n86) );
  CMX2X1 U1608 ( .A0(n710), .A1(C[1]), .S(n18), .Z(n87) );
  CMX2X1 U1609 ( .A0(n652), .A1(C[3]), .S(n18), .Z(n89) );
  CMX2X1 U1610 ( .A0(n654), .A1(C[4]), .S(n18), .Z(n90) );
  CMX2X1 U1611 ( .A0(n656), .A1(C[5]), .S(n18), .Z(n91) );
  CMX2X1 U1612 ( .A0(n226), .A1(C[6]), .S(n18), .Z(n92) );
  CMX2X1 U1613 ( .A0(n227), .A1(C[7]), .S(n18), .Z(n93) );
  CMX2X1 U1614 ( .A0(n225), .A1(C[8]), .S(n18), .Z(n94) );
  CMX2X1 U1615 ( .A0(n362), .A1(C[9]), .S(n18), .Z(n95) );
  CMX2X1 U1616 ( .A0(captC[10]), .A1(C[10]), .S(n18), .Z(n96) );
  CMX2X1 U1617 ( .A0(n511), .A1(C[11]), .S(n18), .Z(n97) );
  CMX2X1 U1618 ( .A0(n658), .A1(C[12]), .S(n18), .Z(n98) );
  CMX2X1 U1619 ( .A0(n661), .A1(C[13]), .S(n18), .Z(n99) );
  CMX2X1 U1620 ( .A0(n650), .A1(C[14]), .S(n18), .Z(n100) );
  CMX2X1 U1621 ( .A0(n664), .A1(C[15]), .S(n18), .Z(n101) );
  CMX2X1 U1622 ( .A0(n667), .A1(C[16]), .S(n18), .Z(n102) );
  CMX2X1 U1623 ( .A0(n670), .A1(C[18]), .S(n18), .Z(n104) );
  CMX2X1 U1624 ( .A0(n673), .A1(C[19]), .S(n18), .Z(n105) );
  CMX2X1 U1625 ( .A0(n676), .A1(C[20]), .S(n18), .Z(n106) );
  CMX2X1 U1626 ( .A0(captC[21]), .A1(C[21]), .S(n18), .Z(n107) );
  CMX2X1 U1627 ( .A0(captC[22]), .A1(C[22]), .S(n18), .Z(n108) );
  CMX2X1 U1628 ( .A0(captC[23]), .A1(C[23]), .S(n18), .Z(n109) );
  CMX2X1 U1629 ( .A0(captC[24]), .A1(C[24]), .S(n18), .Z(n110) );
  CMX2X1 U1630 ( .A0(captC[25]), .A1(C[25]), .S(n18), .Z(n111) );
  CMX2X1 U1631 ( .A0(captC[26]), .A1(C[26]), .S(n18), .Z(n112) );
  CMX2X1 U1632 ( .A0(captC[27]), .A1(C[27]), .S(n18), .Z(n113) );
  CMX2X1 U1633 ( .A0(captC[29]), .A1(C[29]), .S(n18), .Z(n115) );
  CMX2X1 U1634 ( .A0(f27[31]), .A1(f38[31]), .S(rst), .Z(n85) );
  CMX2X1 U1635 ( .A0(f27[30]), .A1(f38[30]), .S(rst), .Z(n84) );
  CMX2X1 U1636 ( .A0(f27[29]), .A1(f38[29]), .S(rst), .Z(n83) );
  CMX2X1 U1637 ( .A0(f27[28]), .A1(f38[28]), .S(rst), .Z(n82) );
  CMX2X1 U1638 ( .A0(f27[27]), .A1(f38[27]), .S(rst), .Z(n81) );
  CMX2X1 U1639 ( .A0(f27[26]), .A1(f38[26]), .S(rst), .Z(n80) );
  CMX2X1 U1640 ( .A0(f27[24]), .A1(f38[24]), .S(rst), .Z(n78) );
  CMX2X1 U1641 ( .A0(f27[23]), .A1(f38[23]), .S(rst), .Z(n77) );
  CMX2X1 U1642 ( .A0(f27[22]), .A1(f38[22]), .S(rst), .Z(n76) );
  CMX2X1 U1643 ( .A0(f27[21]), .A1(f38[21]), .S(rst), .Z(n75) );
  CMX2X1 U1644 ( .A0(f27[20]), .A1(f38[20]), .S(rst), .Z(n74) );
  CMX2X1 U1645 ( .A0(f27[19]), .A1(f38[19]), .S(rst), .Z(n73) );
  CMX2X1 U1646 ( .A0(f27[18]), .A1(f38[18]), .S(rst), .Z(n72) );
  CMX2X1 U1647 ( .A0(f27[17]), .A1(f38[17]), .S(rst), .Z(n71) );
  CMX2X1 U1648 ( .A0(f27[16]), .A1(f38[16]), .S(rst), .Z(n70) );
  CMX2X1 U1649 ( .A0(f27[15]), .A1(f38[15]), .S(rst), .Z(n69) );
  CMX2X1 U1650 ( .A0(f27[14]), .A1(f38[14]), .S(rst), .Z(n68) );
  CMX2X1 U1651 ( .A0(f27[13]), .A1(f38[13]), .S(rst), .Z(n67) );
  CMX2X1 U1652 ( .A0(f27[12]), .A1(f38[12]), .S(rst), .Z(n66) );
  CMX2X1 U1653 ( .A0(f27[11]), .A1(f38[11]), .S(rst), .Z(n65) );
  CMX2X1 U1654 ( .A0(f27[10]), .A1(f38[10]), .S(rst), .Z(n64) );
  CMX2X1 U1655 ( .A0(f27[9]), .A1(f38[9]), .S(rst), .Z(n63) );
  CMX2X1 U1656 ( .A0(f27[8]), .A1(f38[8]), .S(rst), .Z(n62) );
  CMX2X1 U1657 ( .A0(f27[7]), .A1(f38[7]), .S(rst), .Z(n61) );
  CMX2X1 U1658 ( .A0(f27[6]), .A1(f38[6]), .S(rst), .Z(n60) );
  CMX2X1 U1659 ( .A0(f27[5]), .A1(f38[5]), .S(rst), .Z(n59) );
  CMX2X1 U1660 ( .A0(f27[4]), .A1(f38[4]), .S(rst), .Z(n58) );
  CMX2X1 U1661 ( .A0(f27[3]), .A1(f38[3]), .S(rst), .Z(n57) );
  CMX2X1 U1662 ( .A0(f27[2]), .A1(f38[2]), .S(rst), .Z(n56) );
  CMX2X1 U1663 ( .A0(f27[1]), .A1(f38[1]), .S(rst), .Z(n55) );
  CMX2X1 U1664 ( .A0(f27[0]), .A1(f38[0]), .S(rst), .Z(n54) );
  CMX2X1 U1665 ( .A0(s81[5]), .A1(n1406), .S(rst), .Z(n48) );
  CMX2X1 U1666 ( .A0(s81[4]), .A1(n1415), .S(rst), .Z(n49) );
  CMX2X1 U1667 ( .A0(s81[3]), .A1(n1414), .S(rst), .Z(n50) );
  CMX2X1 U1668 ( .A0(s81[2]), .A1(n1413), .S(rst), .Z(n51) );
  CMX2X1 U1669 ( .A0(s81[1]), .A1(n1412), .S(rst), .Z(n52) );
  CMX2X1 U1670 ( .A0(s81[0]), .A1(n1411), .S(rst), .Z(n53) );
  CMX2X1 U1671 ( .A0(s81[6]), .A1(n1407), .S(rst), .Z(n47) );
  CMX2X1 U1672 ( .A0(s81[7]), .A1(n1408), .S(rst), .Z(n46) );
  CMX2X1 U1673 ( .A0(s81[8]), .A1(n1409), .S(rst), .Z(n45) );
  CMX2X1 U1674 ( .A0(s81[9]), .A1(n1410), .S(rst), .Z(n44) );
  CMX2X1 U1675 ( .A0(s81[10]), .A1(n1401), .S(rst), .Z(n43) );
  CMX2X1 U1676 ( .A0(s81[11]), .A1(n1402), .S(rst), .Z(n42) );
  CMX2X1 U1677 ( .A0(s81[12]), .A1(n1403), .S(rst), .Z(n41) );
  CMX2X1 U1678 ( .A0(s81[13]), .A1(n1404), .S(rst), .Z(n40) );
  CMX2X1 U1679 ( .A0(s81[14]), .A1(n1405), .S(rst), .Z(n39) );
  CMX2X1 U1680 ( .A0(s81[15]), .A1(n1396), .S(rst), .Z(n38) );
  CMX2X1 U1681 ( .A0(s81[16]), .A1(n1397), .S(rst), .Z(n37) );
  CMX2X1 U1682 ( .A0(s81[17]), .A1(n1398), .S(rst), .Z(n36) );
  CMX2X1 U1683 ( .A0(s81[18]), .A1(n1399), .S(rst), .Z(n35) );
  CMX2X1 U1684 ( .A0(s81[19]), .A1(n1400), .S(rst), .Z(n34) );
  CMX2X1 U1685 ( .A0(s81[20]), .A1(n1391), .S(rst), .Z(n33) );
  CMX2X1 U1686 ( .A0(s81[21]), .A1(n1392), .S(rst), .Z(n32) );
  CMX2X1 U1687 ( .A0(s81[22]), .A1(n1393), .S(rst), .Z(n31) );
  CMX2X1 U1688 ( .A0(s81[23]), .A1(n1394), .S(rst), .Z(n30) );
  CMX2X1 U1689 ( .A0(s81[24]), .A1(n1395), .S(rst), .Z(n29) );
  CMX2X1 U1690 ( .A0(s81[25]), .A1(n1386), .S(rst), .Z(n28) );
  CMX2X1 U1691 ( .A0(s81[26]), .A1(n1387), .S(rst), .Z(n27) );
  CMX2X1 U1692 ( .A0(s81[27]), .A1(n1388), .S(rst), .Z(n26) );
  CMX2X1 U1693 ( .A0(s81[28]), .A1(n1389), .S(rst), .Z(n25) );
  CMX2X1 U1694 ( .A0(s81[29]), .A1(n1390), .S(rst), .Z(n24) );
  CMX2X1 U1695 ( .A0(s81[30]), .A1(n1384), .S(rst), .Z(n23) );
  CMX2X1 U1696 ( .A0(s81[31]), .A1(n1385), .S(rst), .Z(n22) );
endmodule

